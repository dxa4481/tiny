module tt_um_rebeccargb_universal_decoder (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sg13g2_inv_2 _473_ (.Y(_169_),
    .A(net203));
 sg13g2_inv_1 _474_ (.Y(_180_),
    .A(net226));
 sg13g2_inv_2 _475_ (.Y(_191_),
    .A(net223));
 sg13g2_inv_1 _476_ (.Y(_202_),
    .A(net200));
 sg13g2_inv_2 _477_ (.Y(_212_),
    .A(net199));
 sg13g2_inv_1 _478_ (.Y(_223_),
    .A(net214));
 sg13g2_inv_2 _479_ (.Y(_234_),
    .A(net195));
 sg13g2_nor2_1 _480_ (.A(net204),
    .B(net191),
    .Y(_245_));
 sg13g2_nor2_1 _481_ (.A(net220),
    .B(net217),
    .Y(_255_));
 sg13g2_or2_1 _482_ (.X(_266_),
    .B(net217),
    .A(net221));
 sg13g2_nor2_1 _483_ (.A(net226),
    .B(net223),
    .Y(_277_));
 sg13g2_or2_1 _484_ (.X(_288_),
    .B(net222),
    .A(net225));
 sg13g2_nor2_1 _485_ (.A(net223),
    .B(net2),
    .Y(_298_));
 sg13g2_or2_1 _486_ (.X(_309_),
    .B(net220),
    .A(net224));
 sg13g2_nor4_1 _487_ (.A(net226),
    .B(net223),
    .C(net2),
    .D(net217),
    .Y(_320_));
 sg13g2_nand2_1 _488_ (.Y(_331_),
    .A(_245_),
    .B(net184));
 sg13g2_o21ai_1 _489_ (.B1(net195),
    .Y(_342_),
    .A1(net212),
    .A2(_331_));
 sg13g2_nand2b_2 _490_ (.Y(_352_),
    .B(net207),
    .A_N(net210));
 sg13g2_nand2_2 _491_ (.Y(_363_),
    .A(net203),
    .B(net200));
 sg13g2_and2_1 _492_ (.A(net207),
    .B(net212),
    .X(_374_));
 sg13g2_nand2_2 _493_ (.Y(_384_),
    .A(net207),
    .B(net211));
 sg13g2_nor2_1 _494_ (.A(net210),
    .B(_363_),
    .Y(_395_));
 sg13g2_a22oi_1 _495_ (.Y(_406_),
    .B1(_384_),
    .B2(_395_),
    .A2(_352_),
    .A1(_245_));
 sg13g2_nand2_1 _496_ (.Y(_416_),
    .A(net199),
    .B(_406_));
 sg13g2_a21oi_1 _497_ (.A1(net197),
    .A2(_416_),
    .Y(_425_),
    .B1(net195));
 sg13g2_o21ai_1 _498_ (.B1(_425_),
    .Y(_426_),
    .A1(net198),
    .A2(_416_));
 sg13g2_o21ai_1 _499_ (.B1(_426_),
    .Y(_427_),
    .A1(_212_),
    .A2(_342_));
 sg13g2_nor2b_2 _500_ (.A(net226),
    .B_N(net223),
    .Y(_428_));
 sg13g2_nand2b_2 _501_ (.Y(_429_),
    .B(net222),
    .A_N(net225));
 sg13g2_nor2b_2 _502_ (.A(net220),
    .B_N(net218),
    .Y(_430_));
 sg13g2_nand2b_2 _503_ (.Y(_431_),
    .B(net217),
    .A_N(net221));
 sg13g2_and2_1 _504_ (.A(net219),
    .B(_428_),
    .X(_432_));
 sg13g2_nor2_2 _505_ (.A(net182),
    .B(net180),
    .Y(_433_));
 sg13g2_nand2_1 _506_ (.Y(_434_),
    .A(_428_),
    .B(_430_));
 sg13g2_nand2_1 _507_ (.Y(_435_),
    .A(net219),
    .B(_309_));
 sg13g2_nand4_1 _508_ (.B(net212),
    .C(_309_),
    .A(net219),
    .Y(_436_),
    .D(_434_));
 sg13g2_nand2_1 _509_ (.Y(_437_),
    .A(net190),
    .B(net184));
 sg13g2_nand4_1 _510_ (.B(net196),
    .C(_436_),
    .A(net207),
    .Y(_438_),
    .D(_437_));
 sg13g2_a21oi_1 _511_ (.A1(net199),
    .A2(_331_),
    .Y(_439_),
    .B1(net195));
 sg13g2_nor2_1 _512_ (.A(net193),
    .B(_439_),
    .Y(_440_));
 sg13g2_a22oi_1 _513_ (.Y(_441_),
    .B1(_438_),
    .B2(_440_),
    .A2(_427_),
    .A1(net193));
 sg13g2_inv_1 _514_ (.Y(uo_out[7]),
    .A(_441_));
 sg13g2_and2_1 _515_ (.A(net220),
    .B(net218),
    .X(_442_));
 sg13g2_nand2_1 _516_ (.Y(_443_),
    .A(net221),
    .B(net219));
 sg13g2_nor2_2 _517_ (.A(net183),
    .B(net178),
    .Y(_444_));
 sg13g2_nand2_2 _518_ (.Y(_445_),
    .A(net207),
    .B(net210));
 sg13g2_nand2b_2 _519_ (.Y(_446_),
    .B(net208),
    .A_N(net214));
 sg13g2_inv_1 _520_ (.Y(_447_),
    .A(net177));
 sg13g2_nor2_2 _521_ (.A(net212),
    .B(_445_),
    .Y(_448_));
 sg13g2_nand3b_1 _522_ (.B(net209),
    .C(net208),
    .Y(_449_),
    .A_N(net213));
 sg13g2_nor3_2 _523_ (.A(net182),
    .B(net178),
    .C(net176),
    .Y(_450_));
 sg13g2_nor2_2 _524_ (.A(net189),
    .B(net183),
    .Y(_451_));
 sg13g2_and3_2 _525_ (.X(_452_),
    .A(net208),
    .B(net213),
    .C(net3));
 sg13g2_nand3_1 _526_ (.B(net211),
    .C(net210),
    .A(net207),
    .Y(_453_));
 sg13g2_nor3_1 _527_ (.A(net188),
    .B(net182),
    .C(_453_),
    .Y(_454_));
 sg13g2_o21ai_1 _528_ (.B1(net205),
    .Y(_455_),
    .A1(_450_),
    .A2(_454_));
 sg13g2_nand2b_1 _529_ (.Y(_456_),
    .B(net225),
    .A_N(net222));
 sg13g2_nor2_1 _530_ (.A(net179),
    .B(net174),
    .Y(_457_));
 sg13g2_nor2_2 _531_ (.A(net190),
    .B(_352_),
    .Y(_458_));
 sg13g2_nand3b_1 _532_ (.B(net216),
    .C(net208),
    .Y(_459_),
    .A_N(net209));
 sg13g2_nand2_1 _533_ (.Y(_460_),
    .A(net211),
    .B(net166));
 sg13g2_nor3_2 _534_ (.A(net179),
    .B(net174),
    .C(_459_),
    .Y(_461_));
 sg13g2_nand2b_1 _535_ (.Y(_462_),
    .B(net209),
    .A_N(net208));
 sg13g2_nor2_1 _536_ (.A(net213),
    .B(net173),
    .Y(_463_));
 sg13g2_inv_1 _537_ (.Y(_464_),
    .A(net163));
 sg13g2_nor2_2 _538_ (.A(net224),
    .B(net180),
    .Y(_465_));
 sg13g2_nor2_2 _539_ (.A(net186),
    .B(net181),
    .Y(_466_));
 sg13g2_nand2_1 _540_ (.Y(_467_),
    .A(_277_),
    .B(_430_));
 sg13g2_nor2_2 _541_ (.A(net180),
    .B(net174),
    .Y(_468_));
 sg13g2_and2_1 _542_ (.A(net226),
    .B(net223),
    .X(_469_));
 sg13g2_nand2_2 _543_ (.Y(_470_),
    .A(net225),
    .B(net222));
 sg13g2_nand2b_1 _544_ (.Y(_471_),
    .B(_469_),
    .A_N(net220));
 sg13g2_nor2_2 _545_ (.A(net181),
    .B(net172),
    .Y(_472_));
 sg13g2_or3_1 _546_ (.A(net180),
    .B(_459_),
    .C(net172),
    .X(_000_));
 sg13g2_and4_1 _547_ (.A(net226),
    .B(net222),
    .C(net221),
    .D(net217),
    .X(_001_));
 sg13g2_nand4_1 _548_ (.B(net222),
    .C(net221),
    .A(net225),
    .Y(_002_),
    .D(net217));
 sg13g2_nor2_2 _549_ (.A(net211),
    .B(_352_),
    .Y(_003_));
 sg13g2_nand2_1 _550_ (.Y(_004_),
    .A(net171),
    .B(net159));
 sg13g2_a221oi_1 _551_ (.B2(net165),
    .C1(_461_),
    .B1(_472_),
    .A1(net162),
    .Y(_005_),
    .A2(_465_));
 sg13g2_a21oi_1 _552_ (.A1(_004_),
    .A2(_005_),
    .Y(_006_),
    .B1(net191));
 sg13g2_nand2_1 _553_ (.Y(_007_),
    .A(net161),
    .B(net159));
 sg13g2_nor2_2 _554_ (.A(net187),
    .B(net179),
    .Y(_008_));
 sg13g2_nor3_2 _555_ (.A(net187),
    .B(_384_),
    .C(net178),
    .Y(_009_));
 sg13g2_a22oi_1 _556_ (.Y(_010_),
    .B1(_008_),
    .B2(net165),
    .A2(net159),
    .A1(net161));
 sg13g2_nor3_1 _557_ (.A(net186),
    .B(net181),
    .C(_449_),
    .Y(_011_));
 sg13g2_nor3_1 _558_ (.A(net221),
    .B(net186),
    .C(_449_),
    .Y(_012_));
 sg13g2_a221oi_1 _559_ (.B2(net165),
    .C1(_012_),
    .B1(_008_),
    .A1(net161),
    .Y(_013_),
    .A2(net160));
 sg13g2_nor4_2 _560_ (.A(net211),
    .B(net180),
    .C(net173),
    .Y(_014_),
    .D(net172));
 sg13g2_nor2_1 _561_ (.A(net190),
    .B(net173),
    .Y(_015_));
 sg13g2_nand3b_1 _562_ (.B(net213),
    .C(net209),
    .Y(_016_),
    .A_N(net208));
 sg13g2_nor2b_2 _563_ (.A(net218),
    .B_N(net2),
    .Y(_017_));
 sg13g2_nand2b_2 _564_ (.Y(_018_),
    .B(net221),
    .A_N(net217));
 sg13g2_nor2_1 _565_ (.A(net222),
    .B(net169),
    .Y(_019_));
 sg13g2_nor3_1 _566_ (.A(net224),
    .B(net170),
    .C(net169),
    .Y(_020_));
 sg13g2_nor2_1 _567_ (.A(_014_),
    .B(_020_),
    .Y(_021_));
 sg13g2_nor2_2 _568_ (.A(net189),
    .B(net172),
    .Y(_022_));
 sg13g2_nand3_1 _569_ (.B(net167),
    .C(_022_),
    .A(net205),
    .Y(_023_));
 sg13g2_nor3_2 _570_ (.A(net178),
    .B(net176),
    .C(net174),
    .Y(_024_));
 sg13g2_nand2_1 _571_ (.Y(_025_),
    .A(net205),
    .B(_024_));
 sg13g2_nand3_1 _572_ (.B(net209),
    .C(net166),
    .A(net211),
    .Y(_026_));
 sg13g2_nand2_2 _573_ (.Y(_027_),
    .A(net222),
    .B(net220));
 sg13g2_nor2_2 _574_ (.A(_470_),
    .B(net169),
    .Y(_028_));
 sg13g2_a21oi_1 _575_ (.A1(net163),
    .A2(_028_),
    .Y(_029_),
    .B1(_234_));
 sg13g2_nor3_2 _576_ (.A(net180),
    .B(net177),
    .C(net172),
    .Y(_030_));
 sg13g2_nand2_1 _577_ (.Y(_031_),
    .A(_447_),
    .B(_472_));
 sg13g2_nor4_1 _578_ (.A(net219),
    .B(net209),
    .C(_309_),
    .D(net177),
    .Y(_032_));
 sg13g2_a21oi_1 _579_ (.A1(net171),
    .A2(net157),
    .Y(_033_),
    .B1(_032_));
 sg13g2_nor2_2 _580_ (.A(_429_),
    .B(net168),
    .Y(_034_));
 sg13g2_o21ai_1 _581_ (.B1(net165),
    .Y(_035_),
    .A1(net161),
    .A2(net155));
 sg13g2_nor2_2 _582_ (.A(net175),
    .B(net168),
    .Y(_036_));
 sg13g2_nand3_1 _583_ (.B(net167),
    .C(_036_),
    .A(_363_),
    .Y(_037_));
 sg13g2_o21ai_1 _584_ (.B1(net159),
    .Y(_038_),
    .A1(net155),
    .A2(_036_));
 sg13g2_nor4_1 _585_ (.A(net211),
    .B(net182),
    .C(net180),
    .D(net173),
    .Y(_039_));
 sg13g2_nor3_2 _586_ (.A(_191_),
    .B(net188),
    .C(net170),
    .Y(_040_));
 sg13g2_nor2_1 _587_ (.A(_039_),
    .B(_040_),
    .Y(_041_));
 sg13g2_nor3_2 _588_ (.A(net182),
    .B(_453_),
    .C(net168),
    .Y(_042_));
 sg13g2_nand2_1 _589_ (.Y(_043_),
    .A(_169_),
    .B(_042_));
 sg13g2_nor3_2 _590_ (.A(net176),
    .B(net172),
    .C(net168),
    .Y(_044_));
 sg13g2_nand2b_2 _591_ (.Y(_045_),
    .B(net203),
    .A_N(net200));
 sg13g2_nand3_1 _592_ (.B(net191),
    .C(_044_),
    .A(net203),
    .Y(_046_));
 sg13g2_nor2_2 _593_ (.A(net187),
    .B(net169),
    .Y(_047_));
 sg13g2_nand2_1 _594_ (.Y(_048_),
    .A(_452_),
    .B(_047_));
 sg13g2_nand3_1 _595_ (.B(_452_),
    .C(_047_),
    .A(net203),
    .Y(_049_));
 sg13g2_o21ai_1 _596_ (.B1(_374_),
    .Y(_050_),
    .A1(_468_),
    .A2(_028_));
 sg13g2_o21ai_1 _597_ (.B1(net157),
    .Y(_051_),
    .A1(_465_),
    .A2(net155));
 sg13g2_nor3_1 _598_ (.A(net189),
    .B(_429_),
    .C(net177),
    .Y(_052_));
 sg13g2_nor3_1 _599_ (.A(net186),
    .B(net177),
    .C(net168),
    .Y(_053_));
 sg13g2_nor2_1 _600_ (.A(net188),
    .B(net174),
    .Y(_054_));
 sg13g2_nor3_2 _601_ (.A(net189),
    .B(net176),
    .C(net175),
    .Y(_055_));
 sg13g2_inv_1 _602_ (.Y(_056_),
    .A(_055_));
 sg13g2_nor3_1 _603_ (.A(_052_),
    .B(_053_),
    .C(_055_),
    .Y(_057_));
 sg13g2_nor2_1 _604_ (.A(net206),
    .B(net201),
    .Y(_058_));
 sg13g2_nor2_2 _605_ (.A(_449_),
    .B(_002_),
    .Y(_059_));
 sg13g2_nand2b_1 _606_ (.Y(_060_),
    .B(_059_),
    .A_N(_058_));
 sg13g2_nor3_1 _607_ (.A(net219),
    .B(_309_),
    .C(_384_),
    .Y(_061_));
 sg13g2_a21oi_1 _608_ (.A1(net164),
    .A2(net171),
    .Y(_062_),
    .B1(_061_));
 sg13g2_nor3_2 _609_ (.A(net183),
    .B(net178),
    .C(net170),
    .Y(_063_));
 sg13g2_nor3_2 _610_ (.A(net187),
    .B(net179),
    .C(net170),
    .Y(_064_));
 sg13g2_nor3_2 _611_ (.A(net181),
    .B(_453_),
    .C(net172),
    .Y(_065_));
 sg13g2_nand2_2 _612_ (.Y(_066_),
    .A(_374_),
    .B(_433_));
 sg13g2_nor3_1 _613_ (.A(net188),
    .B(_384_),
    .C(net172),
    .Y(_067_));
 sg13g2_nand2_1 _614_ (.Y(_068_),
    .A(_374_),
    .B(_022_));
 sg13g2_a21oi_1 _615_ (.A1(_066_),
    .A2(_068_),
    .Y(_069_),
    .B1(net200));
 sg13g2_nand3_1 _616_ (.B(net167),
    .C(net155),
    .A(_363_),
    .Y(_070_));
 sg13g2_nand4_1 _617_ (.B(_043_),
    .C(_049_),
    .A(_038_),
    .Y(_071_),
    .D(_070_));
 sg13g2_nand4_1 _618_ (.B(_037_),
    .C(_041_),
    .A(_021_),
    .Y(_072_),
    .D(_062_));
 sg13g2_nand4_1 _619_ (.B(_035_),
    .C(_046_),
    .A(_033_),
    .Y(_073_),
    .D(_050_));
 sg13g2_nand4_1 _620_ (.B(_013_),
    .C(_026_),
    .A(_455_),
    .Y(_074_),
    .D(_057_));
 sg13g2_nor4_1 _621_ (.A(_071_),
    .B(_072_),
    .C(_073_),
    .D(_074_),
    .Y(_075_));
 sg13g2_nand4_1 _622_ (.B(_025_),
    .C(_051_),
    .A(_023_),
    .Y(_076_),
    .D(_060_));
 sg13g2_nor2_1 _623_ (.A(_063_),
    .B(_064_),
    .Y(_077_));
 sg13g2_a21oi_1 _624_ (.A1(net162),
    .A2(net155),
    .Y(_078_),
    .B1(_065_));
 sg13g2_nor3_1 _625_ (.A(net187),
    .B(net180),
    .C(_453_),
    .Y(_079_));
 sg13g2_a221oi_1 _626_ (.B2(_452_),
    .C1(_030_),
    .B1(net161),
    .A1(net166),
    .Y(_080_),
    .A2(net164));
 sg13g2_nand4_1 _627_ (.B(_077_),
    .C(_078_),
    .A(_029_),
    .Y(_081_),
    .D(_080_));
 sg13g2_nor4_1 _628_ (.A(_006_),
    .B(_069_),
    .C(_076_),
    .D(_081_),
    .Y(_082_));
 sg13g2_nor3_2 _629_ (.A(net178),
    .B(_453_),
    .C(net174),
    .Y(_083_));
 sg13g2_a21o_1 _630_ (.A2(net157),
    .A1(net171),
    .B1(_036_),
    .X(_084_));
 sg13g2_nor2_1 _631_ (.A(_047_),
    .B(_063_),
    .Y(_085_));
 sg13g2_a21oi_1 _632_ (.A1(net166),
    .A2(net157),
    .Y(_086_),
    .B1(_022_));
 sg13g2_nand2b_1 _633_ (.Y(_087_),
    .B(_086_),
    .A_N(_084_));
 sg13g2_nor3_1 _634_ (.A(_047_),
    .B(_063_),
    .C(_087_),
    .Y(_088_));
 sg13g2_nand2b_2 _635_ (.Y(_089_),
    .B(net212),
    .A_N(net210));
 sg13g2_nor2_2 _636_ (.A(net207),
    .B(_089_),
    .Y(_090_));
 sg13g2_a21oi_1 _637_ (.A1(net166),
    .A2(net163),
    .Y(_091_),
    .B1(_465_));
 sg13g2_nor2_2 _638_ (.A(_451_),
    .B(_064_),
    .Y(_092_));
 sg13g2_nand2_1 _639_ (.Y(_093_),
    .A(net202),
    .B(_234_));
 sg13g2_nor2_1 _640_ (.A(_083_),
    .B(_093_),
    .Y(_094_));
 sg13g2_nand2_1 _641_ (.Y(_095_),
    .A(_472_),
    .B(_090_));
 sg13g2_nor3_1 _642_ (.A(net155),
    .B(_083_),
    .C(_093_),
    .Y(_096_));
 sg13g2_nand2b_1 _643_ (.Y(_097_),
    .B(_094_),
    .A_N(net155));
 sg13g2_and2_1 _644_ (.A(_095_),
    .B(_096_),
    .X(_098_));
 sg13g2_nor3_1 _645_ (.A(net183),
    .B(net181),
    .C(_453_),
    .Y(_099_));
 sg13g2_nor2_1 _646_ (.A(_450_),
    .B(_099_),
    .Y(_100_));
 sg13g2_nor3_2 _647_ (.A(net187),
    .B(net179),
    .C(net176),
    .Y(_101_));
 sg13g2_nor3_2 _648_ (.A(_384_),
    .B(net182),
    .C(net178),
    .Y(_102_));
 sg13g2_a21oi_1 _649_ (.A1(net210),
    .A2(_030_),
    .Y(_103_),
    .B1(_102_));
 sg13g2_inv_1 _650_ (.Y(_104_),
    .A(_103_));
 sg13g2_a221oi_1 _651_ (.B2(net210),
    .C1(_102_),
    .B1(_030_),
    .A1(_452_),
    .Y(_105_),
    .A2(net171));
 sg13g2_a21oi_1 _652_ (.A1(_432_),
    .A2(_090_),
    .Y(_106_),
    .B1(_039_));
 sg13g2_nand2_1 _653_ (.Y(_107_),
    .A(_105_),
    .B(_106_));
 sg13g2_a21oi_1 _654_ (.A1(_433_),
    .A2(net167),
    .Y(_108_),
    .B1(_014_));
 sg13g2_and2_1 _655_ (.A(_003_),
    .B(_008_),
    .X(_109_));
 sg13g2_o21ai_1 _656_ (.B1(net159),
    .Y(_110_),
    .A1(_472_),
    .A2(_008_));
 sg13g2_nand4_1 _657_ (.B(_092_),
    .C(_108_),
    .A(_091_),
    .Y(_111_),
    .D(_110_));
 sg13g2_nand2b_1 _658_ (.Y(_112_),
    .B(_100_),
    .A_N(_065_));
 sg13g2_nor4_1 _659_ (.A(net224),
    .B(net207),
    .C(net178),
    .D(_089_),
    .Y(_113_));
 sg13g2_nor2_1 _660_ (.A(_101_),
    .B(_113_),
    .Y(_114_));
 sg13g2_a22oi_1 _661_ (.Y(_115_),
    .B1(net159),
    .B2(net166),
    .A2(net165),
    .A1(_433_));
 sg13g2_nand4_1 _662_ (.B(_096_),
    .C(_114_),
    .A(_095_),
    .Y(_116_),
    .D(_115_));
 sg13g2_nor4_1 _663_ (.A(_107_),
    .B(_111_),
    .C(_112_),
    .D(_116_),
    .Y(_117_));
 sg13g2_a22oi_1 _664_ (.Y(_118_),
    .B1(_088_),
    .B2(_117_),
    .A2(_082_),
    .A1(_075_));
 sg13g2_or2_1 _665_ (.X(_119_),
    .B(_118_),
    .A(net194));
 sg13g2_nand2_2 _666_ (.Y(_120_),
    .A(net202),
    .B(net196));
 sg13g2_nand2_1 _667_ (.Y(_121_),
    .A(net212),
    .B(net188));
 sg13g2_or2_1 _668_ (.X(_122_),
    .B(_121_),
    .A(net208));
 sg13g2_a21o_1 _669_ (.A2(net175),
    .A1(net183),
    .B1(net188),
    .X(_123_));
 sg13g2_a21oi_1 _670_ (.A1(net183),
    .A2(net175),
    .Y(_124_),
    .B1(net188));
 sg13g2_mux2_1 _671_ (.A0(net184),
    .A1(net171),
    .S(net190),
    .X(_125_));
 sg13g2_a21oi_1 _672_ (.A1(net214),
    .A2(_124_),
    .Y(_126_),
    .B1(_125_));
 sg13g2_nand2_1 _673_ (.Y(_127_),
    .A(net214),
    .B(_017_));
 sg13g2_a22oi_1 _674_ (.Y(_128_),
    .B1(_469_),
    .B2(_255_),
    .A2(_442_),
    .A1(_428_));
 sg13g2_nand2b_1 _675_ (.Y(_129_),
    .B(net214),
    .A_N(_128_));
 sg13g2_a21o_2 _676_ (.A2(_128_),
    .A1(_467_),
    .B1(net190),
    .X(_130_));
 sg13g2_nor2_2 _677_ (.A(net179),
    .B(_469_),
    .Y(_131_));
 sg13g2_a21oi_1 _678_ (.A1(net224),
    .A2(_430_),
    .Y(_132_),
    .B1(_131_));
 sg13g2_or2_1 _679_ (.X(_133_),
    .B(_132_),
    .A(net215));
 sg13g2_nand4_1 _680_ (.B(_127_),
    .C(_130_),
    .A(_126_),
    .Y(_134_),
    .D(_133_));
 sg13g2_a21oi_1 _681_ (.A1(_122_),
    .A2(_134_),
    .Y(_135_),
    .B1(_120_));
 sg13g2_nor2_1 _682_ (.A(_277_),
    .B(_435_),
    .Y(_136_));
 sg13g2_nand2_1 _683_ (.Y(_137_),
    .A(_234_),
    .B(net6));
 sg13g2_nor3_1 _684_ (.A(_019_),
    .B(_136_),
    .C(_137_),
    .Y(_138_));
 sg13g2_o21ai_1 _685_ (.B1(net193),
    .Y(_139_),
    .A1(_135_),
    .A2(_138_));
 sg13g2_nand3_1 _686_ (.B(_119_),
    .C(_139_),
    .A(net199),
    .Y(_140_));
 sg13g2_xor2_1 _687_ (.B(_140_),
    .A(net197),
    .X(uo_out[6]));
 sg13g2_a221oi_1 _688_ (.B2(net167),
    .C1(_059_),
    .B1(_022_),
    .A1(_451_),
    .Y(_141_),
    .A2(_452_));
 sg13g2_nor2_1 _689_ (.A(net205),
    .B(_141_),
    .Y(_142_));
 sg13g2_nand2_1 _690_ (.Y(_143_),
    .A(net201),
    .B(_064_));
 sg13g2_nand3_1 _691_ (.B(net164),
    .C(net161),
    .A(net192),
    .Y(_144_));
 sg13g2_nand3_1 _692_ (.B(net160),
    .C(_131_),
    .A(net186),
    .Y(_145_));
 sg13g2_a22oi_1 _693_ (.Y(_146_),
    .B1(net156),
    .B2(_447_),
    .A2(net165),
    .A1(_451_));
 sg13g2_nor3_1 _694_ (.A(_180_),
    .B(net217),
    .C(_298_),
    .Y(_147_));
 sg13g2_nand2_1 _695_ (.Y(_148_),
    .A(net160),
    .B(_147_));
 sg13g2_a21oi_1 _696_ (.A1(_001_),
    .A2(net160),
    .Y(_149_),
    .B1(_061_));
 sg13g2_nand4_1 _697_ (.B(_143_),
    .C(_144_),
    .A(_037_),
    .Y(_150_),
    .D(_149_));
 sg13g2_nand3_1 _698_ (.B(_146_),
    .C(_148_),
    .A(_145_),
    .Y(_151_));
 sg13g2_nor3_1 _699_ (.A(_142_),
    .B(_150_),
    .C(_151_),
    .Y(_152_));
 sg13g2_a21oi_2 _700_ (.B1(_052_),
    .Y(_153_),
    .A2(net156),
    .A1(net164));
 sg13g2_nand2_1 _701_ (.Y(_154_),
    .A(net201),
    .B(_065_));
 sg13g2_nor4_1 _702_ (.A(_191_),
    .B(net213),
    .C(net188),
    .D(_462_),
    .Y(_155_));
 sg13g2_nor3_1 _703_ (.A(net225),
    .B(_459_),
    .C(_027_),
    .Y(_156_));
 sg13g2_and3_2 _704_ (.X(_157_),
    .A(net5),
    .B(_469_),
    .C(_017_));
 sg13g2_nor3_1 _705_ (.A(_453_),
    .B(net174),
    .C(net168),
    .Y(_158_));
 sg13g2_nor2_1 _706_ (.A(_450_),
    .B(_158_),
    .Y(_159_));
 sg13g2_nor4_1 _707_ (.A(_450_),
    .B(_024_),
    .C(_042_),
    .D(_158_),
    .Y(_160_));
 sg13g2_nand2_1 _708_ (.Y(_161_),
    .A(_169_),
    .B(_024_));
 sg13g2_nor2_1 _709_ (.A(net205),
    .B(_160_),
    .Y(_162_));
 sg13g2_a221oi_1 _710_ (.B2(net184),
    .C1(_030_),
    .B1(net157),
    .A1(net210),
    .Y(_163_),
    .A2(_009_));
 sg13g2_o21ai_1 _711_ (.B1(net191),
    .Y(_164_),
    .A1(_063_),
    .A2(_083_));
 sg13g2_a22oi_1 _712_ (.Y(_165_),
    .B1(_045_),
    .B2(_101_),
    .A2(_036_),
    .A1(net165));
 sg13g2_nor3_1 _713_ (.A(net219),
    .B(_309_),
    .C(net170),
    .Y(_166_));
 sg13g2_and4_1 _714_ (.A(_049_),
    .B(_163_),
    .C(_164_),
    .D(_165_),
    .X(_167_));
 sg13g2_nor4_2 _715_ (.A(net213),
    .B(net186),
    .C(net173),
    .Y(_168_),
    .D(net169));
 sg13g2_a22oi_1 _716_ (.Y(_170_),
    .B1(_168_),
    .B2(net192),
    .A2(_036_),
    .A1(net164));
 sg13g2_and2_1 _717_ (.A(net196),
    .B(_000_),
    .X(_171_));
 sg13g2_nor4_1 _718_ (.A(_020_),
    .B(_109_),
    .C(_155_),
    .D(_156_),
    .Y(_172_));
 sg13g2_a22oi_1 _719_ (.Y(_173_),
    .B1(_157_),
    .B2(net157),
    .A2(_055_),
    .A1(_169_));
 sg13g2_nor4_1 _720_ (.A(_032_),
    .B(_039_),
    .C(_044_),
    .D(_067_),
    .Y(_174_));
 sg13g2_and2_1 _721_ (.A(_013_),
    .B(_170_),
    .X(_175_));
 sg13g2_and4_1 _722_ (.A(_167_),
    .B(_172_),
    .C(_174_),
    .D(_175_),
    .X(_176_));
 sg13g2_o21ai_1 _723_ (.B1(_154_),
    .Y(_177_),
    .A1(net201),
    .A2(_000_));
 sg13g2_nand4_1 _724_ (.B(_051_),
    .C(_153_),
    .A(_050_),
    .Y(_178_),
    .D(_173_));
 sg13g2_nor3_1 _725_ (.A(_162_),
    .B(_177_),
    .C(_178_),
    .Y(_179_));
 sg13g2_nand4_1 _726_ (.B(_152_),
    .C(_176_),
    .A(net196),
    .Y(_181_),
    .D(_179_));
 sg13g2_a21oi_2 _727_ (.B1(_024_),
    .Y(_182_),
    .A2(_472_),
    .A1(net165));
 sg13g2_inv_1 _728_ (.Y(_183_),
    .A(_182_));
 sg13g2_nor4_1 _729_ (.A(_461_),
    .B(_101_),
    .C(_112_),
    .D(_183_),
    .Y(_184_));
 sg13g2_nor2b_1 _730_ (.A(_009_),
    .B_N(_105_),
    .Y(_185_));
 sg13g2_a221oi_1 _731_ (.B2(_131_),
    .C1(_157_),
    .B1(_090_),
    .A1(_433_),
    .Y(_186_),
    .A2(net158));
 sg13g2_nor4_1 _732_ (.A(_465_),
    .B(_014_),
    .C(net155),
    .D(_084_),
    .Y(_187_));
 sg13g2_a21oi_1 _733_ (.A1(net204),
    .A2(net184),
    .Y(_188_),
    .B1(_093_));
 sg13g2_and4_1 _734_ (.A(_085_),
    .B(_186_),
    .C(_187_),
    .D(_188_),
    .X(_189_));
 sg13g2_nand3_1 _735_ (.B(_185_),
    .C(_189_),
    .A(_184_),
    .Y(_190_));
 sg13g2_a21o_1 _736_ (.A2(_190_),
    .A1(_181_),
    .B1(net194),
    .X(_192_));
 sg13g2_nand2_1 _737_ (.Y(_193_),
    .A(net196),
    .B(_122_));
 sg13g2_nand3_1 _738_ (.B(net216),
    .C(_442_),
    .A(_191_),
    .Y(_194_));
 sg13g2_nand3_1 _739_ (.B(_129_),
    .C(_194_),
    .A(_126_),
    .Y(_195_));
 sg13g2_nor2_1 _740_ (.A(net215),
    .B(_469_),
    .Y(_196_));
 sg13g2_a22oi_1 _741_ (.Y(_197_),
    .B1(_017_),
    .B2(_196_),
    .A2(_430_),
    .A1(net215));
 sg13g2_nor2_1 _742_ (.A(_277_),
    .B(_197_),
    .Y(_198_));
 sg13g2_a22oi_1 _743_ (.Y(_199_),
    .B1(_469_),
    .B2(_017_),
    .A2(_298_),
    .A1(net218));
 sg13g2_a21oi_1 _744_ (.A1(_132_),
    .A2(_199_),
    .Y(_200_),
    .B1(net215));
 sg13g2_nor3_1 _745_ (.A(_195_),
    .B(_198_),
    .C(_200_),
    .Y(_201_));
 sg13g2_nand4_1 _746_ (.B(_445_),
    .C(net177),
    .A(net204),
    .Y(_203_),
    .D(_464_));
 sg13g2_a21oi_1 _747_ (.A1(_169_),
    .A2(net170),
    .Y(_204_),
    .B1(net195));
 sg13g2_nand2_1 _748_ (.Y(_205_),
    .A(net202),
    .B(net193));
 sg13g2_a21oi_1 _749_ (.A1(_203_),
    .A2(_204_),
    .Y(_206_),
    .B1(_205_));
 sg13g2_o21ai_1 _750_ (.B1(_206_),
    .Y(_207_),
    .A1(_193_),
    .A2(_201_));
 sg13g2_nand3_1 _751_ (.B(_192_),
    .C(_207_),
    .A(net199),
    .Y(_208_));
 sg13g2_xor2_1 _752_ (.B(_208_),
    .A(net197),
    .X(uo_out[5]));
 sg13g2_a221oi_1 _753_ (.B2(_451_),
    .C1(_011_),
    .B1(net158),
    .A1(net164),
    .Y(_209_),
    .A2(net161));
 sg13g2_nand2_1 _754_ (.Y(_210_),
    .A(_146_),
    .B(_209_));
 sg13g2_nand2_1 _755_ (.Y(_211_),
    .A(_363_),
    .B(_055_));
 sg13g2_a22oi_1 _756_ (.Y(_213_),
    .B1(_168_),
    .B2(net201),
    .A2(_055_),
    .A1(_363_));
 sg13g2_o21ai_1 _757_ (.B1(net167),
    .Y(_214_),
    .A1(_433_),
    .A2(_028_));
 sg13g2_o21ai_1 _758_ (.B1(_213_),
    .Y(_215_),
    .A1(net203),
    .A2(_214_));
 sg13g2_o21ai_1 _759_ (.B1(_374_),
    .Y(_216_),
    .A1(net184),
    .A2(_028_));
 sg13g2_nand3_1 _760_ (.B(_444_),
    .C(net162),
    .A(net200),
    .Y(_217_));
 sg13g2_nand4_1 _761_ (.B(_171_),
    .C(_216_),
    .A(_153_),
    .Y(_218_),
    .D(_217_));
 sg13g2_a21oi_1 _762_ (.A1(net163),
    .A2(net171),
    .Y(_219_),
    .B1(_454_));
 sg13g2_nand4_1 _763_ (.B(_033_),
    .C(_066_),
    .A(_007_),
    .Y(_220_),
    .D(_219_));
 sg13g2_nor4_1 _764_ (.A(_210_),
    .B(_215_),
    .C(_218_),
    .D(_220_),
    .Y(_221_));
 sg13g2_nand2_1 _765_ (.Y(_222_),
    .A(net225),
    .B(_155_));
 sg13g2_nand2_1 _766_ (.Y(_224_),
    .A(net205),
    .B(_042_));
 sg13g2_nand4_1 _767_ (.B(_159_),
    .C(_222_),
    .A(_025_),
    .Y(_225_),
    .D(_224_));
 sg13g2_a21o_1 _768_ (.A2(net171),
    .A1(net191),
    .B1(_444_),
    .X(_226_));
 sg13g2_a221oi_1 _769_ (.B2(net160),
    .C1(_225_),
    .B1(_226_),
    .A1(_406_),
    .Y(_227_),
    .A2(_059_));
 sg13g2_nor3_1 _770_ (.A(_429_),
    .B(net170),
    .C(net169),
    .Y(_228_));
 sg13g2_o21ai_1 _771_ (.B1(_448_),
    .Y(_229_),
    .A1(_022_),
    .A2(_036_));
 sg13g2_nor4_2 _772_ (.A(net3),
    .B(net183),
    .C(net181),
    .Y(_230_),
    .D(net177));
 sg13g2_nor2_1 _773_ (.A(_228_),
    .B(_230_),
    .Y(_231_));
 sg13g2_a21oi_1 _774_ (.A1(_466_),
    .A2(net158),
    .Y(_232_),
    .B1(_109_));
 sg13g2_a21oi_1 _775_ (.A1(_003_),
    .A2(_147_),
    .Y(_233_),
    .B1(_053_));
 sg13g2_and4_1 _776_ (.A(_229_),
    .B(_231_),
    .C(_232_),
    .D(_233_),
    .X(_235_));
 sg13g2_nand4_1 _777_ (.B(_221_),
    .C(_227_),
    .A(_167_),
    .Y(_236_),
    .D(_235_));
 sg13g2_a21oi_1 _778_ (.A1(net204),
    .A2(net184),
    .Y(_237_),
    .B1(_107_));
 sg13g2_o21ai_1 _779_ (.B1(_092_),
    .Y(_238_),
    .A1(_434_),
    .A2(net170));
 sg13g2_nor4_1 _780_ (.A(net161),
    .B(_009_),
    .C(_097_),
    .D(_238_),
    .Y(_239_));
 sg13g2_nand3_1 _781_ (.B(_237_),
    .C(_239_),
    .A(_184_),
    .Y(_240_));
 sg13g2_nor3_1 _782_ (.A(_444_),
    .B(_468_),
    .C(_047_),
    .Y(_241_));
 sg13g2_or2_1 _783_ (.X(_242_),
    .B(_241_),
    .A(net211));
 sg13g2_nand3_1 _784_ (.B(_130_),
    .C(_242_),
    .A(_460_),
    .Y(_243_));
 sg13g2_a21oi_1 _785_ (.A1(_122_),
    .A2(_243_),
    .Y(_244_),
    .B1(_120_));
 sg13g2_a21oi_1 _786_ (.A1(net226),
    .A2(_027_),
    .Y(_246_),
    .B1(_435_));
 sg13g2_nor3_1 _787_ (.A(_022_),
    .B(_137_),
    .C(_246_),
    .Y(_247_));
 sg13g2_a21o_1 _788_ (.A2(_240_),
    .A1(_236_),
    .B1(net193),
    .X(_248_));
 sg13g2_o21ai_1 _789_ (.B1(net193),
    .Y(_249_),
    .A1(_244_),
    .A2(_247_));
 sg13g2_nand3_1 _790_ (.B(_248_),
    .C(_249_),
    .A(net199),
    .Y(_250_));
 sg13g2_xor2_1 _791_ (.B(_250_),
    .A(net197),
    .X(uo_out[4]));
 sg13g2_a22oi_1 _792_ (.Y(_251_),
    .B1(net157),
    .B2(net166),
    .A2(net162),
    .A1(_444_));
 sg13g2_nor2_1 _793_ (.A(net200),
    .B(_251_),
    .Y(_252_));
 sg13g2_a22oi_1 _794_ (.Y(_253_),
    .B1(_168_),
    .B2(net192),
    .A2(net158),
    .A1(net185));
 sg13g2_a21oi_1 _795_ (.A1(net158),
    .A2(_036_),
    .Y(_254_),
    .B1(_040_));
 sg13g2_nand3_1 _796_ (.B(_253_),
    .C(_254_),
    .A(_154_),
    .Y(_256_));
 sg13g2_nor3_1 _797_ (.A(net181),
    .B(_470_),
    .C(_016_),
    .Y(_257_));
 sg13g2_nand3_1 _798_ (.B(_430_),
    .C(net158),
    .A(net224),
    .Y(_258_));
 sg13g2_nand2_1 _799_ (.Y(_259_),
    .A(net200),
    .B(_083_));
 sg13g2_a21oi_1 _800_ (.A1(_457_),
    .A2(net160),
    .Y(_260_),
    .B1(_158_));
 sg13g2_nand2_1 _801_ (.Y(_261_),
    .A(net163),
    .B(_008_));
 sg13g2_a21oi_1 _802_ (.A1(_446_),
    .A2(_459_),
    .Y(_262_),
    .B1(_002_));
 sg13g2_nand2_1 _803_ (.Y(_263_),
    .A(net162),
    .B(_054_));
 sg13g2_and3_1 _804_ (.X(_264_),
    .A(_050_),
    .B(_066_),
    .C(_263_));
 sg13g2_a21oi_1 _805_ (.A1(_048_),
    .A2(_056_),
    .Y(_265_),
    .B1(_045_));
 sg13g2_nand3_1 _806_ (.B(_468_),
    .C(net157),
    .A(net6),
    .Y(_267_));
 sg13g2_a221oi_1 _807_ (.B2(net184),
    .C1(_262_),
    .B1(net159),
    .A1(net162),
    .Y(_268_),
    .A2(_465_));
 sg13g2_nand3_1 _808_ (.B(_261_),
    .C(_268_),
    .A(_165_),
    .Y(_269_));
 sg13g2_nand3_1 _809_ (.B(_259_),
    .C(_267_),
    .A(_035_),
    .Y(_270_));
 sg13g2_nor4_1 _810_ (.A(_461_),
    .B(_042_),
    .C(_067_),
    .D(_079_),
    .Y(_271_));
 sg13g2_nand3_1 _811_ (.B(_260_),
    .C(_271_),
    .A(_171_),
    .Y(_272_));
 sg13g2_nand4_1 _812_ (.B(_161_),
    .C(_214_),
    .A(_153_),
    .Y(_273_),
    .D(_258_));
 sg13g2_nor4_1 _813_ (.A(_269_),
    .B(_270_),
    .C(_272_),
    .D(_273_),
    .Y(_274_));
 sg13g2_nor3_1 _814_ (.A(_252_),
    .B(_256_),
    .C(_265_),
    .Y(_275_));
 sg13g2_nand4_1 _815_ (.B(_264_),
    .C(_274_),
    .A(_235_),
    .Y(_276_),
    .D(_275_));
 sg13g2_a21oi_1 _816_ (.A1(net206),
    .A2(net185),
    .Y(_278_),
    .B1(_230_));
 sg13g2_a21oi_1 _817_ (.A1(_444_),
    .A2(net163),
    .Y(_279_),
    .B1(_065_));
 sg13g2_nand3_1 _818_ (.B(_182_),
    .C(_279_),
    .A(_110_),
    .Y(_280_));
 sg13g2_a22oi_1 _819_ (.Y(_281_),
    .B1(_090_),
    .B2(net166),
    .A2(_468_),
    .A1(net6));
 sg13g2_nand4_1 _820_ (.B(_106_),
    .C(_278_),
    .A(_095_),
    .Y(_282_),
    .D(_281_));
 sg13g2_nor4_1 _821_ (.A(_087_),
    .B(_104_),
    .C(_280_),
    .D(_282_),
    .Y(_283_));
 sg13g2_nand2_1 _822_ (.Y(_284_),
    .A(_239_),
    .B(_283_));
 sg13g2_a21oi_1 _823_ (.A1(_276_),
    .A2(_284_),
    .Y(_285_),
    .B1(net194));
 sg13g2_nand2_1 _824_ (.Y(_286_),
    .A(_130_),
    .B(_194_));
 sg13g2_o21ai_1 _825_ (.B1(net190),
    .Y(_287_),
    .A1(_022_),
    .A2(_047_));
 sg13g2_nor3_1 _826_ (.A(_223_),
    .B(_451_),
    .C(_028_),
    .Y(_289_));
 sg13g2_a221oi_1 _827_ (.B2(net186),
    .C1(net214),
    .B1(_131_),
    .A1(net218),
    .Y(_290_),
    .A2(_298_));
 sg13g2_o21ai_1 _828_ (.B1(_287_),
    .Y(_291_),
    .A1(_289_),
    .A2(_290_));
 sg13g2_nor2_1 _829_ (.A(_286_),
    .B(_291_),
    .Y(_292_));
 sg13g2_nor2_1 _830_ (.A(_193_),
    .B(_292_),
    .Y(_293_));
 sg13g2_a22oi_1 _831_ (.Y(_294_),
    .B1(net173),
    .B2(net206),
    .A2(net209),
    .A1(net190));
 sg13g2_nor3_1 _832_ (.A(net195),
    .B(net167),
    .C(_294_),
    .Y(_295_));
 sg13g2_nor3_1 _833_ (.A(_205_),
    .B(_293_),
    .C(_295_),
    .Y(_296_));
 sg13g2_nor3_1 _834_ (.A(_212_),
    .B(_285_),
    .C(_296_),
    .Y(_297_));
 sg13g2_xnor2_1 _835_ (.Y(uo_out[3]),
    .A(net197),
    .B(_297_));
 sg13g2_mux2_1 _836_ (.A0(_123_),
    .A1(_199_),
    .S(net190),
    .X(_299_));
 sg13g2_and4_1 _837_ (.A(_130_),
    .B(_194_),
    .C(_287_),
    .D(_299_),
    .X(_300_));
 sg13g2_o21ai_1 _838_ (.B1(net213),
    .Y(_301_),
    .A1(_191_),
    .A2(net169));
 sg13g2_or3_1 _839_ (.A(net213),
    .B(_451_),
    .C(_131_),
    .X(_302_));
 sg13g2_o21ai_1 _840_ (.B1(_302_),
    .Y(_303_),
    .A1(_472_),
    .A2(_301_));
 sg13g2_nand3_1 _841_ (.B(_300_),
    .C(_303_),
    .A(_437_),
    .Y(_304_));
 sg13g2_o21ai_1 _842_ (.B1(_122_),
    .Y(_305_),
    .A1(net206),
    .A2(_437_));
 sg13g2_inv_1 _843_ (.Y(_306_),
    .A(_305_));
 sg13g2_a21oi_1 _844_ (.A1(_304_),
    .A2(_306_),
    .Y(_307_),
    .B1(_120_));
 sg13g2_nand2_1 _845_ (.Y(_308_),
    .A(net219),
    .B(net182));
 sg13g2_o21ai_1 _846_ (.B1(_308_),
    .Y(_310_),
    .A1(_191_),
    .A2(net220));
 sg13g2_a21oi_1 _847_ (.A1(_471_),
    .A2(_310_),
    .Y(_311_),
    .B1(_137_));
 sg13g2_o21ai_1 _848_ (.B1(net8),
    .Y(_312_),
    .A1(_307_),
    .A2(_311_));
 sg13g2_a21o_1 _849_ (.A2(net185),
    .A1(net206),
    .B1(_257_),
    .X(_313_));
 sg13g2_nor4_1 _850_ (.A(_465_),
    .B(_054_),
    .C(_099_),
    .D(_313_),
    .Y(_314_));
 sg13g2_nor2_1 _851_ (.A(_028_),
    .B(_101_),
    .Y(_315_));
 sg13g2_nor2_1 _852_ (.A(_434_),
    .B(net173),
    .Y(_316_));
 sg13g2_nor4_1 _853_ (.A(_028_),
    .B(_065_),
    .C(_101_),
    .D(_316_),
    .Y(_317_));
 sg13g2_nand4_1 _854_ (.B(_098_),
    .C(_314_),
    .A(_088_),
    .Y(_318_),
    .D(_317_));
 sg13g2_o21ai_1 _855_ (.B1(net159),
    .Y(_319_),
    .A1(_028_),
    .A2(_054_));
 sg13g2_nand3_1 _856_ (.B(_214_),
    .C(_319_),
    .A(_050_),
    .Y(_321_));
 sg13g2_nor4_1 _857_ (.A(_011_),
    .B(_228_),
    .C(_230_),
    .D(_257_),
    .Y(_322_));
 sg13g2_nand4_1 _858_ (.B(_021_),
    .C(_031_),
    .A(net196),
    .Y(_323_),
    .D(_322_));
 sg13g2_nor3_1 _859_ (.A(_431_),
    .B(net176),
    .C(net175),
    .Y(_324_));
 sg13g2_nand2_1 _860_ (.Y(_325_),
    .A(net167),
    .B(_468_));
 sg13g2_a21oi_1 _861_ (.A1(net162),
    .A2(_468_),
    .Y(_326_),
    .B1(_166_));
 sg13g2_nand4_1 _862_ (.B(_261_),
    .C(_325_),
    .A(_010_),
    .Y(_327_),
    .D(_326_));
 sg13g2_nor3_1 _863_ (.A(_321_),
    .B(_323_),
    .C(_327_),
    .Y(_328_));
 sg13g2_nand2b_1 _864_ (.Y(_329_),
    .B(_015_),
    .A_N(_199_));
 sg13g2_nand4_1 _865_ (.B(_430_),
    .C(_452_),
    .A(net191),
    .Y(_330_),
    .D(_469_));
 sg13g2_o21ai_1 _866_ (.B1(_330_),
    .Y(_332_),
    .A1(_016_),
    .A2(_199_));
 sg13g2_o21ai_1 _867_ (.B1(_068_),
    .Y(_333_),
    .A1(net203),
    .A2(_048_));
 sg13g2_nand2_1 _868_ (.Y(_334_),
    .A(_468_),
    .B(net160));
 sg13g2_a21oi_1 _869_ (.A1(net204),
    .A2(_101_),
    .Y(_335_),
    .B1(_461_));
 sg13g2_nand2_1 _870_ (.Y(_336_),
    .A(_334_),
    .B(_335_));
 sg13g2_a22oi_1 _871_ (.Y(_337_),
    .B1(_064_),
    .B2(net191),
    .A2(_019_),
    .A1(_458_));
 sg13g2_o21ai_1 _872_ (.B1(net225),
    .Y(_338_),
    .A1(_040_),
    .A2(_061_));
 sg13g2_nand4_1 _873_ (.B(_170_),
    .C(_337_),
    .A(_057_),
    .Y(_339_),
    .D(_338_));
 sg13g2_nor4_1 _874_ (.A(_332_),
    .B(_333_),
    .C(_336_),
    .D(_339_),
    .Y(_340_));
 sg13g2_nand3_1 _875_ (.B(_328_),
    .C(_340_),
    .A(_227_),
    .Y(_341_));
 sg13g2_a21o_1 _876_ (.A2(_341_),
    .A1(_318_),
    .B1(net193),
    .X(_343_));
 sg13g2_nand3_1 _877_ (.B(_312_),
    .C(_343_),
    .A(net199),
    .Y(_344_));
 sg13g2_xor2_1 _878_ (.B(_344_),
    .A(net198),
    .X(uo_out[2]));
 sg13g2_nand3_1 _879_ (.B(net162),
    .C(_468_),
    .A(net191),
    .Y(_345_));
 sg13g2_nand2_1 _880_ (.Y(_346_),
    .A(net200),
    .B(_063_));
 sg13g2_nand3_1 _881_ (.B(_345_),
    .C(_346_),
    .A(_033_),
    .Y(_347_));
 sg13g2_or2_1 _882_ (.X(_348_),
    .B(_059_),
    .A(_011_));
 sg13g2_a221oi_1 _883_ (.B2(_169_),
    .C1(_347_),
    .B1(_348_),
    .A1(net192),
    .Y(_349_),
    .A2(_336_));
 sg13g2_o21ai_1 _884_ (.B1(_259_),
    .Y(_350_),
    .A1(net203),
    .A2(_048_));
 sg13g2_or4_1 _885_ (.A(_053_),
    .B(_155_),
    .C(_156_),
    .D(_230_),
    .X(_351_));
 sg13g2_nand4_1 _886_ (.B(_041_),
    .C(_108_),
    .A(_029_),
    .Y(_353_),
    .D(_145_));
 sg13g2_nor4_1 _887_ (.A(net176),
    .B(net174),
    .C(net168),
    .D(_045_),
    .Y(_354_));
 sg13g2_a221oi_1 _888_ (.B2(_324_),
    .C1(_354_),
    .B1(_058_),
    .A1(net206),
    .Y(_355_),
    .A2(_044_));
 sg13g2_o21ai_1 _889_ (.B1(_355_),
    .Y(_356_),
    .A1(net205),
    .A2(_160_));
 sg13g2_nor4_1 _890_ (.A(_350_),
    .B(_351_),
    .C(_353_),
    .D(_356_),
    .Y(_357_));
 sg13g2_nor4_1 _891_ (.A(_363_),
    .B(net182),
    .C(net176),
    .D(net168),
    .Y(_358_));
 sg13g2_nand2b_1 _892_ (.Y(_359_),
    .B(_337_),
    .A_N(_332_));
 sg13g2_a21oi_1 _893_ (.A1(net158),
    .A2(_047_),
    .Y(_360_),
    .B1(_166_));
 sg13g2_nand4_1 _894_ (.B(_007_),
    .C(_062_),
    .A(_004_),
    .Y(_361_),
    .D(_360_));
 sg13g2_nand4_1 _895_ (.B(_066_),
    .C(_213_),
    .A(_050_),
    .Y(_362_),
    .D(_263_));
 sg13g2_nor4_1 _896_ (.A(_358_),
    .B(_359_),
    .C(_361_),
    .D(_362_),
    .Y(_364_));
 sg13g2_nand3_1 _897_ (.B(_357_),
    .C(_364_),
    .A(_349_),
    .Y(_365_));
 sg13g2_a21oi_1 _898_ (.A1(_008_),
    .A2(_090_),
    .Y(_366_),
    .B1(_450_));
 sg13g2_and4_1 _899_ (.A(_094_),
    .B(_314_),
    .C(_315_),
    .D(_366_),
    .X(_367_));
 sg13g2_nor2_1 _900_ (.A(_014_),
    .B(_238_),
    .Y(_368_));
 sg13g2_nand4_1 _901_ (.B(_086_),
    .C(_367_),
    .A(_085_),
    .Y(_369_),
    .D(_368_));
 sg13g2_a21oi_1 _902_ (.A1(_365_),
    .A2(_369_),
    .Y(_370_),
    .B1(net193));
 sg13g2_a21oi_1 _903_ (.A1(_300_),
    .A2(_303_),
    .Y(_371_),
    .B1(_193_));
 sg13g2_nand3_1 _904_ (.B(net177),
    .C(net173),
    .A(net204),
    .Y(_372_));
 sg13g2_o21ai_1 _905_ (.B1(_372_),
    .Y(_373_),
    .A1(net204),
    .A2(_374_));
 sg13g2_a21oi_1 _906_ (.A1(_089_),
    .A2(_373_),
    .Y(_375_),
    .B1(net195));
 sg13g2_nor3_1 _907_ (.A(_205_),
    .B(_371_),
    .C(_375_),
    .Y(_376_));
 sg13g2_nor3_1 _908_ (.A(_212_),
    .B(_370_),
    .C(_376_),
    .Y(_377_));
 sg13g2_xnor2_1 _909_ (.Y(uo_out[1]),
    .A(net198),
    .B(_377_));
 sg13g2_a21oi_1 _910_ (.A1(_026_),
    .A2(_334_),
    .Y(_378_),
    .B1(net192));
 sg13g2_nor2_1 _911_ (.A(_450_),
    .B(_079_),
    .Y(_379_));
 sg13g2_nor2_1 _912_ (.A(net205),
    .B(_379_),
    .Y(_380_));
 sg13g2_nor4_1 _913_ (.A(_256_),
    .B(_347_),
    .C(_378_),
    .D(_380_),
    .Y(_381_));
 sg13g2_nor3_1 _914_ (.A(_461_),
    .B(_044_),
    .C(_102_),
    .Y(_382_));
 sg13g2_o21ai_1 _915_ (.B1(_433_),
    .Y(_383_),
    .A1(_374_),
    .A2(net163));
 sg13g2_nand4_1 _916_ (.B(_031_),
    .C(_382_),
    .A(net196),
    .Y(_385_),
    .D(_383_));
 sg13g2_nand2b_1 _917_ (.Y(_386_),
    .B(_324_),
    .A_N(_058_));
 sg13g2_o21ai_1 _918_ (.B1(_458_),
    .Y(_387_),
    .A1(_466_),
    .A2(_047_));
 sg13g2_nand2_1 _919_ (.Y(_388_),
    .A(net4),
    .B(_228_));
 sg13g2_nand4_1 _920_ (.B(_386_),
    .C(_387_),
    .A(_329_),
    .Y(_389_),
    .D(_388_));
 sg13g2_nand4_1 _921_ (.B(_211_),
    .C(_224_),
    .A(_182_),
    .Y(_390_),
    .D(_258_));
 sg13g2_nor4_1 _922_ (.A(_333_),
    .B(_385_),
    .C(_389_),
    .D(_390_),
    .Y(_391_));
 sg13g2_nand3_1 _923_ (.B(_381_),
    .C(_391_),
    .A(_152_),
    .Y(_392_));
 sg13g2_nand2_1 _924_ (.Y(_393_),
    .A(net4),
    .B(net156));
 sg13g2_nand4_1 _925_ (.B(_145_),
    .C(_199_),
    .A(_100_),
    .Y(_394_),
    .D(_261_));
 sg13g2_o21ai_1 _926_ (.B1(_393_),
    .Y(_396_),
    .A1(net209),
    .A2(_460_));
 sg13g2_nor4_1 _927_ (.A(_087_),
    .B(_109_),
    .C(_394_),
    .D(_396_),
    .Y(_397_));
 sg13g2_nand4_1 _928_ (.B(_188_),
    .C(_368_),
    .A(_185_),
    .Y(_398_),
    .D(_397_));
 sg13g2_a21o_1 _929_ (.A2(_398_),
    .A1(_392_),
    .B1(net8),
    .X(_399_));
 sg13g2_nor4_1 _930_ (.A(_472_),
    .B(net156),
    .C(_124_),
    .D(_131_),
    .Y(_400_));
 sg13g2_or2_1 _931_ (.X(_401_),
    .B(_400_),
    .A(net214));
 sg13g2_nand3_1 _932_ (.B(net215),
    .C(_430_),
    .A(net224),
    .Y(_402_));
 sg13g2_nand2_1 _933_ (.Y(_403_),
    .A(_127_),
    .B(_402_));
 sg13g2_a22oi_1 _934_ (.Y(_404_),
    .B1(_403_),
    .B2(net186),
    .A2(net185),
    .A1(net214));
 sg13g2_nand3_1 _935_ (.B(_401_),
    .C(_404_),
    .A(_300_),
    .Y(_405_));
 sg13g2_a21oi_1 _936_ (.A1(_122_),
    .A2(_405_),
    .Y(_407_),
    .B1(_120_));
 sg13g2_a21oi_1 _937_ (.A1(net1),
    .A2(net220),
    .Y(_408_),
    .B1(_435_));
 sg13g2_a21oi_1 _938_ (.A1(net223),
    .A2(net169),
    .Y(_409_),
    .B1(_180_));
 sg13g2_nor3_1 _939_ (.A(_137_),
    .B(_408_),
    .C(_409_),
    .Y(_410_));
 sg13g2_o21ai_1 _940_ (.B1(net8),
    .Y(_411_),
    .A1(_407_),
    .A2(_410_));
 sg13g2_nand3_1 _941_ (.B(_399_),
    .C(_411_),
    .A(net199),
    .Y(_412_));
 sg13g2_xor2_1 _942_ (.B(_412_),
    .A(net198),
    .X(uo_out[0]));
 sg13g2_a21oi_1 _943_ (.A1(_245_),
    .A2(_445_),
    .Y(_413_),
    .B1(_212_));
 sg13g2_o21ai_1 _944_ (.B1(_413_),
    .Y(_414_),
    .A1(_363_),
    .A2(_464_));
 sg13g2_xnor2_1 _945_ (.Y(_415_),
    .A(net197),
    .B(_414_));
 sg13g2_nand2_1 _946_ (.Y(_417_),
    .A(net195),
    .B(_121_));
 sg13g2_nand2_1 _947_ (.Y(_418_),
    .A(net194),
    .B(_417_));
 sg13g2_a21oi_1 _948_ (.A1(_234_),
    .A2(_415_),
    .Y(uio_out[1]),
    .B1(_418_));
 sg13g2_nor2_1 _949_ (.A(_442_),
    .B(_121_),
    .Y(_419_));
 sg13g2_o21ai_1 _950_ (.B1(_122_),
    .Y(_420_),
    .A1(_195_),
    .A2(_419_));
 sg13g2_nand2b_1 _951_ (.Y(_421_),
    .B(_420_),
    .A_N(_120_));
 sg13g2_nand4_1 _952_ (.B(net6),
    .C(_027_),
    .A(_234_),
    .Y(_422_),
    .D(_308_));
 sg13g2_nand3_1 _953_ (.B(_421_),
    .C(_422_),
    .A(net7),
    .Y(_423_));
 sg13g2_o21ai_1 _954_ (.B1(net194),
    .Y(_424_),
    .A1(net197),
    .A2(_423_));
 sg13g2_a21oi_1 _955_ (.A1(net197),
    .A2(_423_),
    .Y(uio_out[0]),
    .B1(_424_));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_20 (.L_LO(net20));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _968_ (.A(net194),
    .X(uio_oe[0]));
 sg13g2_buf_1 _969_ (.A(net194),
    .X(uio_oe[1]));
 sg13g2_buf_8 fanout155 (.A(_034_),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(_034_),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net158),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(_015_),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(_003_),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(_466_),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(_463_),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(_458_),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(_457_),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(_448_),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(_018_),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(_018_),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(_016_),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(_001_),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(_470_),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(_462_),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(_456_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_456_),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(_449_),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(_446_),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(_443_),
    .X(net179));
 sg13g2_buf_8 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(_431_),
    .X(net181));
 sg13g2_buf_8 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(_429_),
    .X(net183));
 sg13g2_buf_8 fanout184 (.A(_320_),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(_320_),
    .X(net185));
 sg13g2_buf_8 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_8 fanout187 (.A(_288_),
    .X(net187));
 sg13g2_buf_8 fanout188 (.A(_266_),
    .X(net188));
 sg13g2_buf_1 fanout189 (.A(_266_),
    .X(net189));
 sg13g2_buf_8 fanout190 (.A(_223_),
    .X(net190));
 sg13g2_buf_8 fanout191 (.A(_202_),
    .X(net191));
 sg13g2_buf_1 fanout192 (.A(_202_),
    .X(net192));
 sg13g2_buf_8 fanout193 (.A(net194),
    .X(net193));
 sg13g2_buf_8 fanout194 (.A(net8),
    .X(net194));
 sg13g2_buf_8 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_8 fanout196 (.A(uio_in[6]),
    .X(net196));
 sg13g2_buf_8 fanout197 (.A(uio_in[5]),
    .X(net197));
 sg13g2_buf_1 fanout198 (.A(uio_in[5]),
    .X(net198));
 sg13g2_buf_8 fanout199 (.A(net7),
    .X(net199));
 sg13g2_buf_8 fanout200 (.A(net202),
    .X(net200));
 sg13g2_buf_1 fanout201 (.A(net202),
    .X(net201));
 sg13g2_buf_8 fanout202 (.A(uio_in[3]),
    .X(net202));
 sg13g2_buf_8 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_8 fanout204 (.A(ui_in[7]),
    .X(net204));
 sg13g2_buf_8 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_8 fanout206 (.A(ui_in[7]),
    .X(net206));
 sg13g2_buf_8 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_8 fanout208 (.A(ui_in[6]),
    .X(net208));
 sg13g2_buf_8 fanout209 (.A(net3),
    .X(net209));
 sg13g2_buf_8 fanout210 (.A(net3),
    .X(net210));
 sg13g2_buf_8 fanout211 (.A(ui_in[4]),
    .X(net211));
 sg13g2_buf_8 fanout212 (.A(ui_in[4]),
    .X(net212));
 sg13g2_buf_8 fanout213 (.A(net216),
    .X(net213));
 sg13g2_buf_8 fanout214 (.A(net216),
    .X(net214));
 sg13g2_buf_1 fanout215 (.A(net216),
    .X(net215));
 sg13g2_buf_8 fanout216 (.A(ui_in[4]),
    .X(net216));
 sg13g2_buf_8 fanout217 (.A(ui_in[3]),
    .X(net217));
 sg13g2_buf_1 fanout218 (.A(ui_in[3]),
    .X(net218));
 sg13g2_buf_8 fanout219 (.A(ui_in[3]),
    .X(net219));
 sg13g2_buf_8 fanout220 (.A(net221),
    .X(net220));
 sg13g2_buf_8 fanout221 (.A(net2),
    .X(net221));
 sg13g2_buf_8 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_8 fanout223 (.A(net224),
    .X(net223));
 sg13g2_buf_8 fanout224 (.A(ui_in[1]),
    .X(net224));
 sg13g2_buf_8 fanout225 (.A(net226),
    .X(net225));
 sg13g2_buf_8 fanout226 (.A(net1),
    .X(net226));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[1]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[2]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[4]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_9 (.L_LO(net9));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_decap_4 FILLER_18_156 ();
 sg13g2_fill_2 FILLER_18_160 ();
 sg13g2_decap_4 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_2 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_243 ();
 sg13g2_decap_8 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_4 FILLER_18_283 ();
 sg13g2_decap_4 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_4 FILLER_19_140 ();
 sg13g2_decap_4 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_decap_4 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_178 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_decap_4 FILLER_19_190 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_208 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_decap_4 FILLER_19_252 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_decap_4 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_290 ();
 sg13g2_decap_8 FILLER_19_304 ();
 sg13g2_decap_8 FILLER_19_311 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_8 FILLER_19_332 ();
 sg13g2_decap_4 FILLER_19_339 ();
 sg13g2_fill_2 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_4 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_decap_4 FILLER_20_230 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_decap_8 FILLER_20_262 ();
 sg13g2_decap_4 FILLER_20_269 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_decap_8 FILLER_20_296 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_324 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_4 FILLER_20_360 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_decap_4 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_decap_8 FILLER_21_199 ();
 sg13g2_decap_4 FILLER_21_206 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_decap_4 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_decap_4 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_decap_4 FILLER_21_307 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_2 FILLER_21_321 ();
 sg13g2_fill_2 FILLER_21_331 ();
 sg13g2_fill_1 FILLER_21_333 ();
 sg13g2_fill_2 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_fill_1 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_4 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_4 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_289 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_decap_4 FILLER_22_318 ();
 sg13g2_fill_2 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_343 ();
 sg13g2_fill_2 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_126 ();
 sg13g2_fill_1 FILLER_23_128 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_fill_2 FILLER_23_205 ();
 sg13g2_fill_2 FILLER_23_213 ();
 sg13g2_decap_4 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_decap_4 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_decap_4 FILLER_23_275 ();
 sg13g2_fill_2 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_fill_2 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_fill_2 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_135 ();
 sg13g2_decap_4 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_197 ();
 sg13g2_decap_8 FILLER_24_204 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_decap_4 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_238 ();
 sg13g2_decap_4 FILLER_24_251 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_285 ();
 sg13g2_decap_4 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_318 ();
 sg13g2_decap_4 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_decap_4 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_4 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_fill_2 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_152 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_265 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_decap_8 FILLER_25_276 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_fill_2 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_312 ();
 sg13g2_decap_4 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_decap_4 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_2 FILLER_26_174 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_4 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_decap_4 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_decap_4 FILLER_26_277 ();
 sg13g2_decap_4 FILLER_26_299 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_decap_4 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_355 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_153 ();
 sg13g2_decap_4 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_decap_4 FILLER_27_228 ();
 sg13g2_decap_4 FILLER_27_250 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_fill_2 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_268 ();
 sg13g2_decap_8 FILLER_27_278 ();
 sg13g2_decap_4 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_decap_4 FILLER_27_301 ();
 sg13g2_fill_2 FILLER_27_305 ();
 sg13g2_decap_4 FILLER_27_324 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_353 ();
 sg13g2_fill_2 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_decap_8 FILLER_28_173 ();
 sg13g2_decap_8 FILLER_28_180 ();
 sg13g2_decap_8 FILLER_28_192 ();
 sg13g2_decap_8 FILLER_28_199 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_4 FILLER_28_235 ();
 sg13g2_fill_1 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_268 ();
 sg13g2_decap_8 FILLER_28_275 ();
 sg13g2_fill_1 FILLER_28_291 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_fill_1 FILLER_28_317 ();
 sg13g2_fill_2 FILLER_28_331 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_4 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_137 ();
 sg13g2_decap_4 FILLER_29_155 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_decap_4 FILLER_29_199 ();
 sg13g2_decap_4 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_decap_4 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_decap_4 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_254 ();
 sg13g2_decap_4 FILLER_29_265 ();
 sg13g2_fill_2 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_170 ();
 sg13g2_decap_4 FILLER_30_177 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_4 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_decap_4 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_319 ();
 sg13g2_fill_1 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_fill_2 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_160 ();
 sg13g2_decap_4 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_181 ();
 sg13g2_decap_8 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_206 ();
 sg13g2_fill_1 FILLER_31_208 ();
 sg13g2_decap_8 FILLER_31_236 ();
 sg13g2_decap_4 FILLER_31_243 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_299 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_fill_2 FILLER_31_346 ();
 sg13g2_decap_4 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_393 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_4 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_149 ();
 sg13g2_decap_4 FILLER_32_156 ();
 sg13g2_decap_4 FILLER_32_179 ();
 sg13g2_fill_2 FILLER_32_183 ();
 sg13g2_decap_8 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_221 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_240 ();
 sg13g2_decap_8 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_267 ();
 sg13g2_decap_8 FILLER_32_275 ();
 sg13g2_decap_8 FILLER_32_282 ();
 sg13g2_decap_4 FILLER_32_289 ();
 sg13g2_decap_4 FILLER_32_319 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_378 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_4 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_144 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_decap_4 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_194 ();
 sg13g2_decap_4 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_decap_4 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_decap_8 FILLER_33_269 ();
 sg13g2_fill_1 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_decap_4 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_decap_4 FILLER_33_344 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_decap_4 FILLER_33_358 ();
 sg13g2_fill_2 FILLER_33_362 ();
 sg13g2_decap_4 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_4 FILLER_34_178 ();
 sg13g2_decap_4 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_fill_2 FILLER_34_208 ();
 sg13g2_fill_1 FILLER_34_210 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_227 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_decap_4 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_348 ();
 sg13g2_decap_4 FILLER_34_377 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_decap_4 FILLER_34_387 ();
 sg13g2_fill_2 FILLER_34_391 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_4 FILLER_35_161 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_decap_4 FILLER_35_200 ();
 sg13g2_fill_1 FILLER_35_204 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_decap_4 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_8 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_decap_4 FILLER_35_333 ();
 sg13g2_fill_2 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_350 ();
 sg13g2_decap_4 FILLER_35_372 ();
 sg13g2_fill_2 FILLER_35_376 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_fill_2 FILLER_36_207 ();
 sg13g2_fill_1 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_216 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_fill_2 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_247 ();
 sg13g2_decap_4 FILLER_36_254 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_293 ();
 sg13g2_decap_4 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_349 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_4 FILLER_36_390 ();
 sg13g2_fill_2 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_decap_4 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_250 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_decap_8 FILLER_37_293 ();
 sg13g2_decap_8 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_307 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_100 ();
 sg13g2_decap_8 FILLER_38_107 ();
 sg13g2_decap_4 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_118 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_171 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_4 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_238 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_4 FILLER_38_347 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
endmodule
