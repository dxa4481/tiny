module tt_um_chip_rom (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire \addr_counter[0] ;
 wire \addr_counter[1] ;
 wire \addr_counter[2] ;
 wire \addr_counter[3] ;
 wire \addr_counter[4] ;
 wire \addr_counter[5] ;
 wire \addr_counter[6] ;
 wire \addr_counter[7] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire clknet_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net17;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net61;
 wire net62;
 wire net63;
 wire net64;

 sg13g2_inv_4 _193_ (.A(net60),
    .Y(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _194_ (.VDD(VPWR),
    .Y(_137_),
    .A(net39),
    .VSS(VGND));
 sg13g2_inv_1 _195_ (.VDD(VPWR),
    .Y(_000_),
    .A(net33),
    .VSS(VGND));
 sg13g2_and2_1 _196_ (.A(net58),
    .B(net4),
    .X(_138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _197_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net56),
    .A2(\addr_counter[3] ),
    .Y(_139_),
    .B1(_138_));
 sg13g2_mux2_1 _198_ (.A0(\addr_counter[3] ),
    .A1(net4),
    .S(net58),
    .X(_140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _199_ (.A0(\addr_counter[2] ),
    .A1(net3),
    .S(net59),
    .X(_141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _200_ (.Y(_142_),
    .A(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _201_ (.A(net52),
    .B(net48),
    .Y(_143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _202_ (.A(net58),
    .B(net6),
    .X(_144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _203_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_144_),
    .Y(_145_),
    .A2(\addr_counter[5] ),
    .A1(net56));
 sg13g2_a21o_2 _204_ (.A2(\addr_counter[5] ),
    .A1(net56),
    .B1(_144_),
    .X(_146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _205_ (.A(_143_),
    .B(_145_),
    .Y(_147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _206_ (.A(net57),
    .B(net7),
    .X(_148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _207_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_148_),
    .Y(_149_),
    .A2(\addr_counter[6] ),
    .A1(net56));
 sg13g2_a21o_2 _208_ (.A2(\addr_counter[6] ),
    .A1(net56),
    .B1(_148_),
    .X(_150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _209_ (.A(net57),
    .B(net5),
    .X(_151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _210_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_151_),
    .Y(_152_),
    .A2(\addr_counter[4] ),
    .A1(net56));
 sg13g2_a21o_2 _211_ (.A2(\addr_counter[4] ),
    .A1(net56),
    .B1(_151_),
    .X(_153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _212_ (.A(_145_),
    .B(_152_),
    .Y(_154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _213_ (.Y(_155_),
    .A(net47),
    .B(_153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _214_ (.Y(_156_),
    .A(net46),
    .B(_155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _215_ (.A(_147_),
    .B(_156_),
    .Y(_157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _216_ (.A(net57),
    .B(net1),
    .X(_158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _217_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_158_),
    .Y(_159_),
    .A2(\addr_counter[0] ),
    .A1(_008_));
 sg13g2_mux2_1 _218_ (.A0(\addr_counter[0] ),
    .A1(net1),
    .S(net57),
    .X(_160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _219_ (.A(net50),
    .B(net43),
    .Y(_161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _220_ (.Y(_162_),
    .A(net54),
    .B(_159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _221_ (.Y(_163_),
    .A(net45),
    .B(_162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _222_ (.A(net57),
    .B(\addr_counter[1] ),
    .Y(_164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _223_ (.A(net2),
    .B_N(net57),
    .Y(_165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _224_ (.A0(\addr_counter[1] ),
    .A1(net2),
    .S(net57),
    .X(_166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _225_ (.A(net43),
    .B_N(net41),
    .Y(_167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _226_ (.B(net41),
    .A(net43),
    .X(_168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _227_ (.A(net49),
    .B_N(net41),
    .Y(_169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _228_ (.A(net49),
    .B_N(net43),
    .Y(_170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _229_ (.A(net54),
    .B(_168_),
    .C(_169_),
    .Y(_171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _230_ (.Y(_172_),
    .A(net49),
    .B(_168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _231_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net43),
    .C1(net45),
    .B1(_169_),
    .A1(_142_),
    .Y(_173_),
    .A2(_161_));
 sg13g2_o21ai_1 _232_ (.B1(_173_),
    .VDD(VPWR),
    .Y(_174_),
    .VSS(VGND),
    .A1(_161_),
    .A2(_172_));
 sg13g2_o21ai_1 _233_ (.B1(_174_),
    .VDD(VPWR),
    .Y(_175_),
    .VSS(VGND),
    .A1(_163_),
    .A2(_171_));
 sg13g2_nor2_2 _234_ (.A(net50),
    .B(_170_),
    .Y(_176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _235_ (.A(net41),
    .B_N(net49),
    .Y(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _236_ (.Y(_178_),
    .A(net49),
    .B(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _237_ (.A(net48),
    .B(net42),
    .Y(_179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _238_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_180_),
    .B(net42),
    .A(net48));
 sg13g2_xor2_1 _239_ (.B(net41),
    .A(_141_),
    .X(_181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _240_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_182_),
    .B(_181_),
    .A(net44));
 sg13g2_nand2_2 _241_ (.Y(_183_),
    .A(net49),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _242_ (.A(_181_),
    .B_N(_183_),
    .Y(_184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _243_ (.Y(_185_),
    .B(_183_),
    .A_N(_181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _244_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_186_),
    .B(net44),
    .A(net48));
 sg13g2_nor2b_2 _245_ (.A(net44),
    .B_N(net48),
    .Y(_187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _246_ (.Y(_188_),
    .A(_159_),
    .B(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _247_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_159_),
    .A2(_177_),
    .Y(_189_),
    .B1(net55));
 sg13g2_a221oi_1 _248_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_189_),
    .C1(net45),
    .B1(_186_),
    .A1(_176_),
    .Y(_190_),
    .A2(_185_));
 sg13g2_nor3_1 _249_ (.A(net50),
    .B(_170_),
    .C(_177_),
    .Y(_191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _250_ (.Y(_192_),
    .B(net45),
    .A_N(_191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _251_ (.Y(_016_),
    .A(net43),
    .B(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _252_ (.B(net44),
    .C(net42),
    .A(net48),
    .Y(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _253_ (.A(net48),
    .B(net44),
    .C(_164_),
    .D(_165_),
    .X(_018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _254_ (.Y(_019_),
    .A(_017_),
    .B(_018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _255_ (.B1(net47),
    .VDD(VPWR),
    .Y(_020_),
    .VSS(VGND),
    .A1(_192_),
    .A2(_019_));
 sg13g2_nor2_2 _256_ (.A(_146_),
    .B(_153_),
    .Y(_021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _257_ (.Y(_022_),
    .A(_145_),
    .B(_152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _258_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net52),
    .A2(_187_),
    .Y(_023_),
    .B1(_022_));
 sg13g2_nand2b_1 _259_ (.Y(_024_),
    .B(_023_),
    .A_N(_143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _260_ (.B1(_024_),
    .VDD(VPWR),
    .Y(_025_),
    .VSS(VGND),
    .A1(_190_),
    .A2(_020_));
 sg13g2_a22oi_1 _261_ (.Y(_026_),
    .B1(_025_),
    .B2(_149_),
    .A2(_175_),
    .A1(_157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _262_ (.A(net57),
    .B(net8),
    .X(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _263_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_027_),
    .Y(_028_),
    .A2(\addr_counter[7] ),
    .A1(net56));
 sg13g2_inv_1 _264_ (.VDD(VPWR),
    .Y(_029_),
    .A(_028_),
    .VSS(VGND));
 sg13g2_nor2_2 _265_ (.A(_155_),
    .B(_028_),
    .Y(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _266_ (.A(net53),
    .B(net44),
    .C(_181_),
    .D(_030_),
    .X(_031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _267_ (.A0(_028_),
    .A1(_031_),
    .S(_026_),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _268_ (.A(net54),
    .B(_179_),
    .C(_187_),
    .Y(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _269_ (.B(_030_),
    .C(_032_),
    .A(net46),
    .Y(_033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _270_ (.Y(_034_),
    .A(net53),
    .B(_018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _271_ (.B(_017_),
    .C(_018_),
    .A(net52),
    .Y(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _272_ (.A(net52),
    .B(_179_),
    .Y(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _273_ (.Y(_037_),
    .A(net55),
    .B(_180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _274_ (.B1(_035_),
    .VDD(VPWR),
    .Y(_038_),
    .VSS(VGND),
    .A1(_167_),
    .A2(_037_));
 sg13g2_nand2_1 _275_ (.Y(_039_),
    .A(_021_),
    .B(_038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _276_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_036_),
    .C1(_155_),
    .B1(_188_),
    .A1(net52),
    .Y(_040_),
    .A2(_182_));
 sg13g2_nor2_2 _277_ (.A(_145_),
    .B(_153_),
    .Y(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _278_ (.Y(_042_),
    .A(net47),
    .B(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _279_ (.A(net54),
    .B(_172_),
    .Y(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _280_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_161_),
    .A2(_179_),
    .Y(_044_),
    .B1(_043_));
 sg13g2_o21ai_1 _281_ (.B1(_039_),
    .VDD(VPWR),
    .Y(_045_),
    .VSS(VGND),
    .A1(_042_),
    .A2(_044_));
 sg13g2_nor3_1 _282_ (.A(net46),
    .B(_040_),
    .C(_045_),
    .Y(_046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _283_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_188_),
    .A2(_036_),
    .Y(_047_),
    .B1(_043_));
 sg13g2_nor2_2 _284_ (.A(net47),
    .B(net45),
    .Y(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _285_ (.A(_047_),
    .B_N(_048_),
    .Y(_049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _286_ (.B1(_188_),
    .VDD(VPWR),
    .Y(_050_),
    .VSS(VGND),
    .A1(_161_),
    .A2(_036_));
 sg13g2_nand3_1 _287_ (.B(_034_),
    .C(_050_),
    .A(_021_),
    .Y(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _288_ (.B(_177_),
    .C(_041_),
    .A(net54),
    .Y(_052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _289_ (.B(_051_),
    .C(_052_),
    .A(_150_),
    .Y(_053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _290_ (.B1(_028_),
    .VDD(VPWR),
    .Y(_054_),
    .VSS(VGND),
    .A1(_049_),
    .A2(_053_));
 sg13g2_o21ai_1 _291_ (.B1(_033_),
    .VDD(VPWR),
    .Y(net10),
    .VSS(VGND),
    .A1(_046_),
    .A2(_054_));
 sg13g2_nand3_1 _292_ (.B(net46),
    .C(_030_),
    .A(net53),
    .Y(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _293_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_056_),
    .B(_055_),
    .A(_185_));
 sg13g2_nand4_1 _294_ (.B(_180_),
    .C(_017_),
    .A(net52),
    .Y(_057_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_018_));
 sg13g2_and2_1 _295_ (.A(net55),
    .B(_186_),
    .X(_058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _296_ (.Y(_059_),
    .A(net42),
    .B(_058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _297_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_057_),
    .A2(_059_),
    .Y(_060_),
    .B1(_022_));
 sg13g2_nand2_1 _298_ (.Y(_061_),
    .A(_161_),
    .B(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _299_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_159_),
    .A2(_177_),
    .Y(_062_),
    .B1(_170_));
 sg13g2_nor2_1 _300_ (.A(net50),
    .B(_169_),
    .Y(_063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _301_ (.B1(_062_),
    .VDD(VPWR),
    .Y(_064_),
    .VSS(VGND),
    .A1(net50),
    .A2(_168_));
 sg13g2_a21oi_1 _302_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_061_),
    .A2(_064_),
    .Y(_065_),
    .B1(_155_));
 sg13g2_nand2_1 _303_ (.Y(_066_),
    .A(net51),
    .B(_184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _304_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_037_),
    .A2(_066_),
    .Y(_067_),
    .B1(_042_));
 sg13g2_nor4_1 _305_ (.A(net46),
    .B(_060_),
    .C(_065_),
    .D(_067_),
    .Y(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _306_ (.B1(net46),
    .VDD(VPWR),
    .Y(_069_),
    .VSS(VGND),
    .A1(_153_),
    .A2(_061_));
 sg13g2_nor2_1 _307_ (.A(_161_),
    .B(_168_),
    .Y(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _308_ (.A(net45),
    .B(_170_),
    .C(_070_),
    .Y(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _309_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net50),
    .C1(_163_),
    .B1(_181_),
    .A1(net43),
    .Y(_072_),
    .A2(_179_));
 sg13g2_nor3_1 _310_ (.A(net47),
    .B(_071_),
    .C(_072_),
    .Y(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _311_ (.B1(_028_),
    .VDD(VPWR),
    .Y(_074_),
    .VSS(VGND),
    .A1(_069_),
    .A2(_073_));
 sg13g2_o21ai_1 _312_ (.B1(_056_),
    .VDD(VPWR),
    .Y(net11),
    .VSS(VGND),
    .A1(_068_),
    .A2(_074_));
 sg13g2_nor2_2 _313_ (.A(net42),
    .B(_187_),
    .Y(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _314_ (.A(net54),
    .B(net49),
    .Y(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _315_ (.Y(_077_),
    .A(net50),
    .B(_142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _316_ (.B1(_077_),
    .VDD(VPWR),
    .Y(_078_),
    .VSS(VGND),
    .A1(_162_),
    .A2(_178_));
 sg13g2_o21ai_1 _317_ (.B1(_021_),
    .VDD(VPWR),
    .Y(_079_),
    .VSS(VGND),
    .A1(_075_),
    .A2(_078_));
 sg13g2_nor3_1 _318_ (.A(net51),
    .B(_159_),
    .C(_169_),
    .Y(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _319_ (.A(net50),
    .B(_169_),
    .X(_081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _320_ (.B1(_041_),
    .VDD(VPWR),
    .Y(_082_),
    .VSS(VGND),
    .A1(_080_),
    .A2(_081_));
 sg13g2_nand2b_1 _321_ (.Y(_083_),
    .B(_176_),
    .A_N(_167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _322_ (.A2(_083_),
    .A1(_066_),
    .B1(_155_),
    .X(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _323_ (.B(_079_),
    .C(_082_),
    .A(_149_),
    .Y(_085_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_084_));
 sg13g2_and4_1 _324_ (.A(net51),
    .B(_178_),
    .C(_183_),
    .D(_016_),
    .X(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _325_ (.B1(_048_),
    .VDD(VPWR),
    .Y(_087_),
    .VSS(VGND),
    .A1(_080_),
    .A2(_086_));
 sg13g2_nor2_1 _326_ (.A(net54),
    .B(_167_),
    .Y(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _327_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_183_),
    .A2(_088_),
    .Y(_089_),
    .B1(net47));
 sg13g2_nand2b_1 _328_ (.Y(_090_),
    .B(_089_),
    .A_N(_192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _329_ (.B(_041_),
    .C(_075_),
    .A(_176_),
    .Y(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _330_ (.B(_087_),
    .C(_090_),
    .A(net46),
    .Y(_092_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_091_));
 sg13g2_nand3_1 _331_ (.B(_085_),
    .C(_092_),
    .A(_028_),
    .Y(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _332_ (.B1(_093_),
    .VDD(VPWR),
    .Y(net12),
    .VSS(VGND),
    .A1(_184_),
    .A2(_055_));
 sg13g2_xnor2_1 _333_ (.Y(_094_),
    .A(_142_),
    .B(_168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _334_ (.Y(_095_),
    .A(_037_),
    .B(_094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _335_ (.Y(_096_),
    .B(_032_),
    .A_N(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _336_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_168_),
    .A2(_063_),
    .Y(_097_),
    .B1(_042_));
 sg13g2_a221oi_1 _337_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_097_),
    .C1(_023_),
    .B1(_096_),
    .A1(_154_),
    .Y(_098_),
    .A2(_095_));
 sg13g2_nor2_1 _338_ (.A(_150_),
    .B(_098_),
    .Y(_099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _339_ (.B1(_143_),
    .VDD(VPWR),
    .Y(_100_),
    .VSS(VGND),
    .A1(_159_),
    .A2(net42));
 sg13g2_nand2_1 _340_ (.Y(_101_),
    .A(_057_),
    .B(_100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _341_ (.B1(_189_),
    .VDD(VPWR),
    .Y(_102_),
    .VSS(VGND),
    .A1(net48),
    .A2(_168_));
 sg13g2_a21oi_1 _342_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_172_),
    .A2(_058_),
    .Y(_103_),
    .B1(_153_));
 sg13g2_a221oi_1 _343_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_103_),
    .C1(net47),
    .B1(_102_),
    .A1(_153_),
    .Y(_104_),
    .A2(_101_));
 sg13g2_nor2b_1 _344_ (.A(_104_),
    .B_N(_157_),
    .Y(_105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _345_ (.B1(_028_),
    .VDD(VPWR),
    .Y(_106_),
    .VSS(VGND),
    .A1(_099_),
    .A2(_105_));
 sg13g2_o21ai_1 _346_ (.B1(_106_),
    .VDD(VPWR),
    .Y(net13),
    .VSS(VGND),
    .A1(_177_),
    .A2(_055_));
 sg13g2_nand2_1 _347_ (.Y(_107_),
    .A(net55),
    .B(_182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _348_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_034_),
    .A2(_107_),
    .Y(_108_),
    .B1(_145_));
 sg13g2_or2_1 _349_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_109_),
    .B(_183_),
    .A(net41));
 sg13g2_a21o_1 _350_ (.A2(_109_),
    .A1(net55),
    .B1(_032_),
    .X(_110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _351_ (.A2(_110_),
    .A1(_152_),
    .B1(_108_),
    .X(_111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _352_ (.B(_178_),
    .C(_183_),
    .A(net54),
    .Y(_112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _353_ (.Y(_113_),
    .A(net47),
    .B(_112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _354_ (.A(net52),
    .B(net45),
    .C(_109_),
    .Y(_114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _355_ (.A(_156_),
    .B(_114_),
    .Y(_115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _356_ (.Y(_116_),
    .B1(_113_),
    .B2(_115_),
    .A2(_111_),
    .A1(_149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _357_ (.B(_183_),
    .C(net42),
    .Y(_117_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_055_));
 sg13g2_o21ai_1 _358_ (.B1(_117_),
    .VDD(VPWR),
    .Y(net14),
    .VSS(VGND),
    .A1(_029_),
    .A2(_116_));
 sg13g2_a21oi_1 _359_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_162_),
    .A2(_016_),
    .Y(_118_),
    .B1(_169_));
 sg13g2_o21ai_1 _360_ (.B1(_048_),
    .VDD(VPWR),
    .Y(_119_),
    .VSS(VGND),
    .A1(_076_),
    .A2(_118_));
 sg13g2_nand2_1 _361_ (.Y(_120_),
    .A(net51),
    .B(_109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _362_ (.B(_037_),
    .C(_120_),
    .A(_162_),
    .Y(_121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _363_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_021_),
    .A2(_121_),
    .Y(_122_),
    .B1(_069_));
 sg13g2_o21ai_1 _364_ (.B1(_041_),
    .VDD(VPWR),
    .Y(_123_),
    .VSS(VGND),
    .A1(net52),
    .A2(_017_));
 sg13g2_nor2_1 _365_ (.A(_043_),
    .B(_123_),
    .Y(_124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _366_ (.Y(_125_),
    .A(_016_),
    .B(_077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _367_ (.B1(_021_),
    .VDD(VPWR),
    .Y(_126_),
    .VSS(VGND),
    .A1(_063_),
    .A2(_125_));
 sg13g2_a21oi_1 _368_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_176_),
    .A2(_075_),
    .Y(_127_),
    .B1(_155_));
 sg13g2_nor3_1 _369_ (.A(net46),
    .B(_124_),
    .C(_127_),
    .Y(_128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _370_ (.Y(_129_),
    .B1(_126_),
    .B2(_128_),
    .A2(_122_),
    .A1(_119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _371_ (.A(_030_),
    .B(_086_),
    .X(_130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _372_ (.A0(_130_),
    .A1(_028_),
    .S(_129_),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _373_ (.A(_055_),
    .B(_075_),
    .Y(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _374_ (.B(net36),
    .A(net33),
    .X(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _375_ (.B(net33),
    .C(net36),
    .A(net63),
    .Y(_131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _376_ (.A2(net36),
    .A1(net33),
    .B1(net63),
    .X(_132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _377_ (.A(_131_),
    .B(_132_),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _378_ (.A(_137_),
    .B(_131_),
    .Y(_133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _379_ (.Y(_003_),
    .A(net39),
    .B(_131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _380_ (.A(net37),
    .B(_133_),
    .X(_134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _381_ (.B(_133_),
    .A(net37),
    .X(_004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _382_ (.B(_134_),
    .A(net61),
    .X(_005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _383_ (.B(net64),
    .C(_134_),
    .A(net61),
    .Y(_135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _384_ (.A2(_134_),
    .A1(net61),
    .B1(net64),
    .X(_136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _385_ (.A(_135_),
    .B(_136_),
    .X(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _386_ (.Y(_007_),
    .A(net34),
    .B(_135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _387_ (.VDD(VPWR),
    .Y(_009_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _388_ (.VDD(VPWR),
    .Y(_010_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _389_ (.VDD(VPWR),
    .Y(_011_),
    .A(net60),
    .VSS(VGND));
 sg13g2_inv_1 _390_ (.VDD(VPWR),
    .Y(_012_),
    .A(net60),
    .VSS(VGND));
 sg13g2_inv_1 _391_ (.VDD(VPWR),
    .Y(_013_),
    .A(net60),
    .VSS(VGND));
 sg13g2_inv_1 _392_ (.VDD(VPWR),
    .Y(_014_),
    .A(net60),
    .VSS(VGND));
 sg13g2_inv_1 _393_ (.VDD(VPWR),
    .Y(_015_),
    .A(net60),
    .VSS(VGND));
 sg13g2_dfrbpq_2 _394_ (.RESET_B(_008_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_000_),
    .Q(\addr_counter[0] ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _395_ (.RESET_B(_009_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_001_),
    .Q(\addr_counter[1] ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _396_ (.RESET_B(_010_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_002_),
    .Q(\addr_counter[2] ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _397_ (.RESET_B(_011_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net40),
    .Q(\addr_counter[3] ),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _398_ (.RESET_B(_012_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net38),
    .Q(\addr_counter[4] ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _399_ (.RESET_B(_013_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net62),
    .Q(\addr_counter[5] ),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _400_ (.RESET_B(_014_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_006_),
    .Q(\addr_counter[6] ),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _401_ (.RESET_B(_015_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net35),
    .Q(\addr_counter[7] ),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_tielo tt_um_chip_rom_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net18));
 sg13g2_tielo tt_um_chip_rom_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net19));
 sg13g2_tielo tt_um_chip_rom_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net20));
 sg13g2_tielo tt_um_chip_rom_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net21));
 sg13g2_tielo tt_um_chip_rom_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net22));
 sg13g2_tielo tt_um_chip_rom_23 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net23));
 sg13g2_tielo tt_um_chip_rom_24 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net24));
 sg13g2_tielo tt_um_chip_rom_25 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net25));
 sg13g2_tielo tt_um_chip_rom_26 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net26));
 sg13g2_tielo tt_um_chip_rom_27 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net27));
 sg13g2_tielo tt_um_chip_rom_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net28));
 sg13g2_tielo tt_um_chip_rom_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net29));
 sg13g2_tielo tt_um_chip_rom_30 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net30));
 sg13g2_tielo tt_um_chip_rom_31 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net31));
 sg13g2_tielo tt_um_chip_rom_32 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net32));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout41 (.A(_166_),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout42 (.A(_166_),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout43 (.A(_160_),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout44 (.A(_160_),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout45 (.A(_152_),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout46 (.A(_150_),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout47 (.A(_146_),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout48 (.A(_141_),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout49 (.A(_141_),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout50 (.A(net53),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout51 (.A(net53),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout52 (.A(net53),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout53 (.A(_140_),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout54 (.A(_139_),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout55 (.A(_139_),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout56 (.A(_008_),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout57 (.A(net58),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout58 (.A(net59),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout59 (.A(net60),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout60 (.A(rst_n),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo tt_um_chip_rom_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net17));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload0 (.A(clknet_1_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\addr_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold2 (.A(\addr_counter[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold3 (.A(_007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold4 (.A(\addr_counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold5 (.A(\addr_counter[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold6 (.A(_004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold7 (.A(\addr_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold8 (.A(_003_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold9 (.A(\addr_counter[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold10 (.A(_005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold11 (.A(\addr_counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold12 (.A(\addr_counter[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_407 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule
