module tt_mux (k_one,
    k_zero,
    addr,
    spine_iw,
    spine_ow,
    um_ena,
    um_iw,
    um_k_zero,
    um_ow,
    um_pg_ena);
 output k_one;
 output k_zero;
 input [3:0] addr;
 input [29:0] spine_iw;
 output [25:0] spine_ow;
 output [11:0] um_ena;
 output [215:0] um_iw;
 output [11:0] um_k_zero;
 input [287:0] um_ow;
 output [11:0] um_pg_ena;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire \block[0].genblk1.grp_sel_buf_I.a ;
 wire \block[0].genblk1.grp_sel_buf_I.z ;
 wire \block[0].genblk1.l_tbe ;
 wire \block[0].genblk1.mux4_I[0].x ;
 wire \block[0].genblk1.mux4_I[10].x ;
 wire \block[0].genblk1.mux4_I[11].x ;
 wire \block[0].genblk1.mux4_I[12].x ;
 wire \block[0].genblk1.mux4_I[13].x ;
 wire \block[0].genblk1.mux4_I[14].x ;
 wire \block[0].genblk1.mux4_I[15].x ;
 wire \block[0].genblk1.mux4_I[16].x ;
 wire \block[0].genblk1.mux4_I[17].x ;
 wire \block[0].genblk1.mux4_I[18].x ;
 wire \block[0].genblk1.mux4_I[19].x ;
 wire \block[0].genblk1.mux4_I[1].x ;
 wire \block[0].genblk1.mux4_I[20].x ;
 wire \block[0].genblk1.mux4_I[21].x ;
 wire \block[0].genblk1.mux4_I[22].x ;
 wire \block[0].genblk1.mux4_I[23].x ;
 wire \block[0].genblk1.mux4_I[2].x ;
 wire \block[0].genblk1.mux4_I[3].x ;
 wire \block[0].genblk1.mux4_I[4].x ;
 wire \block[0].genblk1.mux4_I[5].x ;
 wire \block[0].genblk1.mux4_I[6].x ;
 wire \block[0].genblk1.mux4_I[7].x ;
 wire \block[0].genblk1.mux4_I[8].x ;
 wire \block[0].genblk1.mux4_I[9].x ;
 wire \block[0].genblk1.mux4_sel_buf_I[0].a ;
 wire \block[0].genblk1.mux4_sel_buf_I[0].z ;
 wire \block[0].genblk1.mux4_sel_buf_I[1].a ;
 wire \block[0].genblk1.mux4_sel_buf_I[1].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[0].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[10].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[11].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[12].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[13].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[14].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[15].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[16].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[17].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[18].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[19].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[1].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[20].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[21].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[22].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[23].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[2].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[3].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[4].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[5].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[6].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[7].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[8].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[9].z ;
 wire \block[0].l_ena ;
 wire \block[0].l_ena_0_I.a ;
 wire \block[0].tie_I.lo ;
 wire \block[0].zbuf_ena_I.z ;
 wire \block[0].zbuf_iw_I[0].a ;
 wire \block[0].zbuf_iw_I[0].z ;
 wire \block[0].zbuf_iw_I[10].a ;
 wire \block[0].zbuf_iw_I[10].z ;
 wire \block[0].zbuf_iw_I[11].a ;
 wire \block[0].zbuf_iw_I[11].z ;
 wire \block[0].zbuf_iw_I[12].a ;
 wire \block[0].zbuf_iw_I[12].z ;
 wire \block[0].zbuf_iw_I[13].a ;
 wire \block[0].zbuf_iw_I[13].z ;
 wire \block[0].zbuf_iw_I[14].a ;
 wire \block[0].zbuf_iw_I[14].z ;
 wire \block[0].zbuf_iw_I[15].a ;
 wire \block[0].zbuf_iw_I[15].z ;
 wire \block[0].zbuf_iw_I[16].a ;
 wire \block[0].zbuf_iw_I[16].z ;
 wire \block[0].zbuf_iw_I[17].a ;
 wire \block[0].zbuf_iw_I[17].z ;
 wire \block[0].zbuf_iw_I[1].a ;
 wire \block[0].zbuf_iw_I[1].z ;
 wire \block[0].zbuf_iw_I[2].a ;
 wire \block[0].zbuf_iw_I[2].z ;
 wire \block[0].zbuf_iw_I[3].a ;
 wire \block[0].zbuf_iw_I[3].z ;
 wire \block[0].zbuf_iw_I[4].a ;
 wire \block[0].zbuf_iw_I[4].z ;
 wire \block[0].zbuf_iw_I[5].a ;
 wire \block[0].zbuf_iw_I[5].z ;
 wire \block[0].zbuf_iw_I[6].a ;
 wire \block[0].zbuf_iw_I[6].z ;
 wire \block[0].zbuf_iw_I[7].a ;
 wire \block[0].zbuf_iw_I[7].z ;
 wire \block[0].zbuf_iw_I[8].a ;
 wire \block[0].zbuf_iw_I[8].z ;
 wire \block[0].zbuf_iw_I[9].a ;
 wire \block[0].zbuf_iw_I[9].z ;
 wire \block[0].zbuf_pg_ena_I.z ;
 wire \block[10].l_ena ;
 wire \block[10].l_ena_0_I.a ;
 wire \block[10].tie_I.lo ;
 wire \block[10].zbuf_ena_I.z ;
 wire \block[10].zbuf_iw_I[0].z ;
 wire \block[10].zbuf_iw_I[10].z ;
 wire \block[10].zbuf_iw_I[11].z ;
 wire \block[10].zbuf_iw_I[12].z ;
 wire \block[10].zbuf_iw_I[13].z ;
 wire \block[10].zbuf_iw_I[14].z ;
 wire \block[10].zbuf_iw_I[15].z ;
 wire \block[10].zbuf_iw_I[16].z ;
 wire \block[10].zbuf_iw_I[17].z ;
 wire \block[10].zbuf_iw_I[1].z ;
 wire \block[10].zbuf_iw_I[2].z ;
 wire \block[10].zbuf_iw_I[3].z ;
 wire \block[10].zbuf_iw_I[4].z ;
 wire \block[10].zbuf_iw_I[5].z ;
 wire \block[10].zbuf_iw_I[6].z ;
 wire \block[10].zbuf_iw_I[7].z ;
 wire \block[10].zbuf_iw_I[8].z ;
 wire \block[10].zbuf_iw_I[9].z ;
 wire \block[10].zbuf_pg_ena_I.z ;
 wire \block[11].l_ena ;
 wire \block[11].l_ena_0_I.a ;
 wire \block[11].tie_I.lo ;
 wire \block[11].zbuf_ena_I.z ;
 wire \block[11].zbuf_iw_I[0].z ;
 wire \block[11].zbuf_iw_I[10].z ;
 wire \block[11].zbuf_iw_I[11].z ;
 wire \block[11].zbuf_iw_I[12].z ;
 wire \block[11].zbuf_iw_I[13].z ;
 wire \block[11].zbuf_iw_I[14].z ;
 wire \block[11].zbuf_iw_I[15].z ;
 wire \block[11].zbuf_iw_I[16].z ;
 wire \block[11].zbuf_iw_I[17].z ;
 wire \block[11].zbuf_iw_I[1].z ;
 wire \block[11].zbuf_iw_I[2].z ;
 wire \block[11].zbuf_iw_I[3].z ;
 wire \block[11].zbuf_iw_I[4].z ;
 wire \block[11].zbuf_iw_I[5].z ;
 wire \block[11].zbuf_iw_I[6].z ;
 wire \block[11].zbuf_iw_I[7].z ;
 wire \block[11].zbuf_iw_I[8].z ;
 wire \block[11].zbuf_iw_I[9].z ;
 wire \block[11].zbuf_pg_ena_I.z ;
 wire \block[1].l_ena ;
 wire \block[1].l_ena_0_I.a ;
 wire \block[1].tie_I.lo ;
 wire \block[1].zbuf_ena_I.z ;
 wire \block[1].zbuf_iw_I[0].z ;
 wire \block[1].zbuf_iw_I[10].z ;
 wire \block[1].zbuf_iw_I[11].z ;
 wire \block[1].zbuf_iw_I[12].z ;
 wire \block[1].zbuf_iw_I[13].z ;
 wire \block[1].zbuf_iw_I[14].z ;
 wire \block[1].zbuf_iw_I[15].z ;
 wire \block[1].zbuf_iw_I[16].z ;
 wire \block[1].zbuf_iw_I[17].z ;
 wire \block[1].zbuf_iw_I[1].z ;
 wire \block[1].zbuf_iw_I[2].z ;
 wire \block[1].zbuf_iw_I[3].z ;
 wire \block[1].zbuf_iw_I[4].z ;
 wire \block[1].zbuf_iw_I[5].z ;
 wire \block[1].zbuf_iw_I[6].z ;
 wire \block[1].zbuf_iw_I[7].z ;
 wire \block[1].zbuf_iw_I[8].z ;
 wire \block[1].zbuf_iw_I[9].z ;
 wire \block[1].zbuf_pg_ena_I.z ;
 wire \block[2].l_ena ;
 wire \block[2].l_ena_0_I.a ;
 wire \block[2].tie_I.lo ;
 wire \block[2].zbuf_ena_I.z ;
 wire \block[2].zbuf_iw_I[0].z ;
 wire \block[2].zbuf_iw_I[10].z ;
 wire \block[2].zbuf_iw_I[11].z ;
 wire \block[2].zbuf_iw_I[12].z ;
 wire \block[2].zbuf_iw_I[13].z ;
 wire \block[2].zbuf_iw_I[14].z ;
 wire \block[2].zbuf_iw_I[15].z ;
 wire \block[2].zbuf_iw_I[16].z ;
 wire \block[2].zbuf_iw_I[17].z ;
 wire \block[2].zbuf_iw_I[1].z ;
 wire \block[2].zbuf_iw_I[2].z ;
 wire \block[2].zbuf_iw_I[3].z ;
 wire \block[2].zbuf_iw_I[4].z ;
 wire \block[2].zbuf_iw_I[5].z ;
 wire \block[2].zbuf_iw_I[6].z ;
 wire \block[2].zbuf_iw_I[7].z ;
 wire \block[2].zbuf_iw_I[8].z ;
 wire \block[2].zbuf_iw_I[9].z ;
 wire \block[2].zbuf_pg_ena_I.z ;
 wire \block[3].l_ena ;
 wire \block[3].l_ena_0_I.a ;
 wire \block[3].tie_I.lo ;
 wire \block[3].zbuf_ena_I.z ;
 wire \block[3].zbuf_iw_I[0].z ;
 wire \block[3].zbuf_iw_I[10].z ;
 wire \block[3].zbuf_iw_I[11].z ;
 wire \block[3].zbuf_iw_I[12].z ;
 wire \block[3].zbuf_iw_I[13].z ;
 wire \block[3].zbuf_iw_I[14].z ;
 wire \block[3].zbuf_iw_I[15].z ;
 wire \block[3].zbuf_iw_I[16].z ;
 wire \block[3].zbuf_iw_I[17].z ;
 wire \block[3].zbuf_iw_I[1].z ;
 wire \block[3].zbuf_iw_I[2].z ;
 wire \block[3].zbuf_iw_I[3].z ;
 wire \block[3].zbuf_iw_I[4].z ;
 wire \block[3].zbuf_iw_I[5].z ;
 wire \block[3].zbuf_iw_I[6].z ;
 wire \block[3].zbuf_iw_I[7].z ;
 wire \block[3].zbuf_iw_I[8].z ;
 wire \block[3].zbuf_iw_I[9].z ;
 wire \block[3].zbuf_pg_ena_I.z ;
 wire \block[4].genblk1.grp_sel_buf_I.a ;
 wire \block[4].genblk1.grp_sel_buf_I.z ;
 wire \block[4].genblk1.l_tbe ;
 wire \block[4].genblk1.mux4_I[0].x ;
 wire \block[4].genblk1.mux4_I[10].x ;
 wire \block[4].genblk1.mux4_I[11].x ;
 wire \block[4].genblk1.mux4_I[12].x ;
 wire \block[4].genblk1.mux4_I[13].x ;
 wire \block[4].genblk1.mux4_I[14].x ;
 wire \block[4].genblk1.mux4_I[15].x ;
 wire \block[4].genblk1.mux4_I[16].x ;
 wire \block[4].genblk1.mux4_I[17].x ;
 wire \block[4].genblk1.mux4_I[18].x ;
 wire \block[4].genblk1.mux4_I[19].x ;
 wire \block[4].genblk1.mux4_I[1].x ;
 wire \block[4].genblk1.mux4_I[20].x ;
 wire \block[4].genblk1.mux4_I[21].x ;
 wire \block[4].genblk1.mux4_I[22].x ;
 wire \block[4].genblk1.mux4_I[23].x ;
 wire \block[4].genblk1.mux4_I[2].x ;
 wire \block[4].genblk1.mux4_I[3].x ;
 wire \block[4].genblk1.mux4_I[4].x ;
 wire \block[4].genblk1.mux4_I[5].x ;
 wire \block[4].genblk1.mux4_I[6].x ;
 wire \block[4].genblk1.mux4_I[7].x ;
 wire \block[4].genblk1.mux4_I[8].x ;
 wire \block[4].genblk1.mux4_I[9].x ;
 wire \block[4].genblk1.mux4_sel_buf_I[0].z ;
 wire \block[4].genblk1.mux4_sel_buf_I[1].z ;
 wire \block[4].l_ena ;
 wire \block[4].l_ena_0_I.a ;
 wire \block[4].tie_I.lo ;
 wire \block[4].zbuf_ena_I.z ;
 wire \block[4].zbuf_iw_I[0].z ;
 wire \block[4].zbuf_iw_I[10].z ;
 wire \block[4].zbuf_iw_I[11].z ;
 wire \block[4].zbuf_iw_I[12].z ;
 wire \block[4].zbuf_iw_I[13].z ;
 wire \block[4].zbuf_iw_I[14].z ;
 wire \block[4].zbuf_iw_I[15].z ;
 wire \block[4].zbuf_iw_I[16].z ;
 wire \block[4].zbuf_iw_I[17].z ;
 wire \block[4].zbuf_iw_I[1].z ;
 wire \block[4].zbuf_iw_I[2].z ;
 wire \block[4].zbuf_iw_I[3].z ;
 wire \block[4].zbuf_iw_I[4].z ;
 wire \block[4].zbuf_iw_I[5].z ;
 wire \block[4].zbuf_iw_I[6].z ;
 wire \block[4].zbuf_iw_I[7].z ;
 wire \block[4].zbuf_iw_I[8].z ;
 wire \block[4].zbuf_iw_I[9].z ;
 wire \block[4].zbuf_pg_ena_I.z ;
 wire \block[5].l_ena ;
 wire \block[5].l_ena_0_I.a ;
 wire \block[5].tie_I.lo ;
 wire \block[5].zbuf_ena_I.z ;
 wire \block[5].zbuf_iw_I[0].z ;
 wire \block[5].zbuf_iw_I[10].z ;
 wire \block[5].zbuf_iw_I[11].z ;
 wire \block[5].zbuf_iw_I[12].z ;
 wire \block[5].zbuf_iw_I[13].z ;
 wire \block[5].zbuf_iw_I[14].z ;
 wire \block[5].zbuf_iw_I[15].z ;
 wire \block[5].zbuf_iw_I[16].z ;
 wire \block[5].zbuf_iw_I[17].z ;
 wire \block[5].zbuf_iw_I[1].z ;
 wire \block[5].zbuf_iw_I[2].z ;
 wire \block[5].zbuf_iw_I[3].z ;
 wire \block[5].zbuf_iw_I[4].z ;
 wire \block[5].zbuf_iw_I[5].z ;
 wire \block[5].zbuf_iw_I[6].z ;
 wire \block[5].zbuf_iw_I[7].z ;
 wire \block[5].zbuf_iw_I[8].z ;
 wire \block[5].zbuf_iw_I[9].z ;
 wire \block[5].zbuf_pg_ena_I.z ;
 wire \block[6].l_ena ;
 wire \block[6].l_ena_0_I.a ;
 wire \block[6].tie_I.lo ;
 wire \block[6].zbuf_ena_I.z ;
 wire \block[6].zbuf_iw_I[0].z ;
 wire \block[6].zbuf_iw_I[10].z ;
 wire \block[6].zbuf_iw_I[11].z ;
 wire \block[6].zbuf_iw_I[12].z ;
 wire \block[6].zbuf_iw_I[13].z ;
 wire \block[6].zbuf_iw_I[14].z ;
 wire \block[6].zbuf_iw_I[15].z ;
 wire \block[6].zbuf_iw_I[16].z ;
 wire \block[6].zbuf_iw_I[17].z ;
 wire \block[6].zbuf_iw_I[1].z ;
 wire \block[6].zbuf_iw_I[2].z ;
 wire \block[6].zbuf_iw_I[3].z ;
 wire \block[6].zbuf_iw_I[4].z ;
 wire \block[6].zbuf_iw_I[5].z ;
 wire \block[6].zbuf_iw_I[6].z ;
 wire \block[6].zbuf_iw_I[7].z ;
 wire \block[6].zbuf_iw_I[8].z ;
 wire \block[6].zbuf_iw_I[9].z ;
 wire \block[6].zbuf_pg_ena_I.z ;
 wire \block[7].l_ena ;
 wire \block[7].l_ena_0_I.a ;
 wire \block[7].tie_I.lo ;
 wire \block[7].zbuf_ena_I.z ;
 wire \block[7].zbuf_iw_I[0].z ;
 wire \block[7].zbuf_iw_I[10].z ;
 wire \block[7].zbuf_iw_I[11].z ;
 wire \block[7].zbuf_iw_I[12].z ;
 wire \block[7].zbuf_iw_I[13].z ;
 wire \block[7].zbuf_iw_I[14].z ;
 wire \block[7].zbuf_iw_I[15].z ;
 wire \block[7].zbuf_iw_I[16].z ;
 wire \block[7].zbuf_iw_I[17].z ;
 wire \block[7].zbuf_iw_I[1].z ;
 wire \block[7].zbuf_iw_I[2].z ;
 wire \block[7].zbuf_iw_I[3].z ;
 wire \block[7].zbuf_iw_I[4].z ;
 wire \block[7].zbuf_iw_I[5].z ;
 wire \block[7].zbuf_iw_I[6].z ;
 wire \block[7].zbuf_iw_I[7].z ;
 wire \block[7].zbuf_iw_I[8].z ;
 wire \block[7].zbuf_iw_I[9].z ;
 wire \block[7].zbuf_pg_ena_I.z ;
 wire \block[8].genblk1.grp_sel_buf_I.a ;
 wire \block[8].genblk1.grp_sel_buf_I.z ;
 wire \block[8].genblk1.l_tbe ;
 wire \block[8].genblk1.mux4_I[0].x ;
 wire \block[8].genblk1.mux4_I[10].x ;
 wire \block[8].genblk1.mux4_I[11].x ;
 wire \block[8].genblk1.mux4_I[12].x ;
 wire \block[8].genblk1.mux4_I[13].x ;
 wire \block[8].genblk1.mux4_I[14].x ;
 wire \block[8].genblk1.mux4_I[15].x ;
 wire \block[8].genblk1.mux4_I[16].x ;
 wire \block[8].genblk1.mux4_I[17].x ;
 wire \block[8].genblk1.mux4_I[18].x ;
 wire \block[8].genblk1.mux4_I[19].x ;
 wire \block[8].genblk1.mux4_I[1].x ;
 wire \block[8].genblk1.mux4_I[20].x ;
 wire \block[8].genblk1.mux4_I[21].x ;
 wire \block[8].genblk1.mux4_I[22].x ;
 wire \block[8].genblk1.mux4_I[23].x ;
 wire \block[8].genblk1.mux4_I[2].x ;
 wire \block[8].genblk1.mux4_I[3].x ;
 wire \block[8].genblk1.mux4_I[4].x ;
 wire \block[8].genblk1.mux4_I[5].x ;
 wire \block[8].genblk1.mux4_I[6].x ;
 wire \block[8].genblk1.mux4_I[7].x ;
 wire \block[8].genblk1.mux4_I[8].x ;
 wire \block[8].genblk1.mux4_I[9].x ;
 wire \block[8].genblk1.mux4_sel_buf_I[0].z ;
 wire \block[8].genblk1.mux4_sel_buf_I[1].z ;
 wire \block[8].l_ena ;
 wire \block[8].l_ena_0_I.a ;
 wire \block[8].tie_I.lo ;
 wire \block[8].zbuf_ena_I.z ;
 wire \block[8].zbuf_iw_I[0].z ;
 wire \block[8].zbuf_iw_I[10].z ;
 wire \block[8].zbuf_iw_I[11].z ;
 wire \block[8].zbuf_iw_I[12].z ;
 wire \block[8].zbuf_iw_I[13].z ;
 wire \block[8].zbuf_iw_I[14].z ;
 wire \block[8].zbuf_iw_I[15].z ;
 wire \block[8].zbuf_iw_I[16].z ;
 wire \block[8].zbuf_iw_I[17].z ;
 wire \block[8].zbuf_iw_I[1].z ;
 wire \block[8].zbuf_iw_I[2].z ;
 wire \block[8].zbuf_iw_I[3].z ;
 wire \block[8].zbuf_iw_I[4].z ;
 wire \block[8].zbuf_iw_I[5].z ;
 wire \block[8].zbuf_iw_I[6].z ;
 wire \block[8].zbuf_iw_I[7].z ;
 wire \block[8].zbuf_iw_I[8].z ;
 wire \block[8].zbuf_iw_I[9].z ;
 wire \block[8].zbuf_pg_ena_I.z ;
 wire \block[9].l_ena ;
 wire \block[9].l_ena_0_I.a ;
 wire \block[9].tie_I.lo ;
 wire \block[9].zbuf_ena_I.z ;
 wire \block[9].zbuf_iw_I[0].z ;
 wire \block[9].zbuf_iw_I[10].z ;
 wire \block[9].zbuf_iw_I[11].z ;
 wire \block[9].zbuf_iw_I[12].z ;
 wire \block[9].zbuf_iw_I[13].z ;
 wire \block[9].zbuf_iw_I[14].z ;
 wire \block[9].zbuf_iw_I[15].z ;
 wire \block[9].zbuf_iw_I[16].z ;
 wire \block[9].zbuf_iw_I[17].z ;
 wire \block[9].zbuf_iw_I[1].z ;
 wire \block[9].zbuf_iw_I[2].z ;
 wire \block[9].zbuf_iw_I[3].z ;
 wire \block[9].zbuf_iw_I[4].z ;
 wire \block[9].zbuf_iw_I[5].z ;
 wire \block[9].zbuf_iw_I[6].z ;
 wire \block[9].zbuf_iw_I[7].z ;
 wire \block[9].zbuf_iw_I[8].z ;
 wire \block[9].zbuf_iw_I[9].z ;
 wire \block[9].zbuf_pg_ena_I.z ;
 wire \branch_addr_match_buf_I[0].z ;
 wire \branch_addr_match_buf_I[1].z ;
 wire \branch_addr_match_buf_I[2].z ;
 wire \branch_addr_match_buf_I[3].z ;
 wire \branch_ena_buf_I.z ;
 wire branch_sel;
 wire \branch_sel_buf_I.a ;
 wire branch_sel_n;
 wire branch_sel_n_tbe;
 wire branch_sel_tbe;
 wire \buf_bus_ena_I.z ;
 wire \buf_bus_sel_I[2].z ;
 wire \buf_bus_sel_I[3].z ;
 wire \buf_bus_sel_I[4].z ;
 wire \buf_spine_ow_I[0].z ;
 wire \buf_spine_ow_I[10].z ;
 wire \buf_spine_ow_I[11].z ;
 wire \buf_spine_ow_I[12].z ;
 wire \buf_spine_ow_I[13].z ;
 wire \buf_spine_ow_I[14].z ;
 wire \buf_spine_ow_I[15].z ;
 wire \buf_spine_ow_I[16].z ;
 wire \buf_spine_ow_I[17].z ;
 wire \buf_spine_ow_I[18].z ;
 wire \buf_spine_ow_I[19].z ;
 wire \buf_spine_ow_I[1].z ;
 wire \buf_spine_ow_I[20].z ;
 wire \buf_spine_ow_I[21].z ;
 wire \buf_spine_ow_I[22].z ;
 wire \buf_spine_ow_I[23].z ;
 wire \buf_spine_ow_I[2].z ;
 wire \buf_spine_ow_I[3].z ;
 wire \buf_spine_ow_I[4].z ;
 wire \buf_spine_ow_I[5].z ;
 wire \buf_spine_ow_I[6].z ;
 wire \buf_spine_ow_I[7].z ;
 wire \buf_spine_ow_I[8].z ;
 wire \buf_spine_ow_I[9].z ;
 wire \bus_pull_ow_I[0].a ;
 wire so_gh;
 wire so_gl;
 wire \tbuf_spine_ow_I[0].z ;
 wire \tbuf_spine_ow_I[10].z ;
 wire \tbuf_spine_ow_I[11].z ;
 wire \tbuf_spine_ow_I[12].z ;
 wire \tbuf_spine_ow_I[13].z ;
 wire \tbuf_spine_ow_I[14].z ;
 wire \tbuf_spine_ow_I[15].z ;
 wire \tbuf_spine_ow_I[16].z ;
 wire \tbuf_spine_ow_I[17].z ;
 wire \tbuf_spine_ow_I[18].z ;
 wire \tbuf_spine_ow_I[19].z ;
 wire \tbuf_spine_ow_I[1].z ;
 wire \tbuf_spine_ow_I[20].z ;
 wire \tbuf_spine_ow_I[21].z ;
 wire \tbuf_spine_ow_I[22].z ;
 wire \tbuf_spine_ow_I[23].z ;
 wire \tbuf_spine_ow_I[2].z ;
 wire \tbuf_spine_ow_I[3].z ;
 wire \tbuf_spine_ow_I[4].z ;
 wire \tbuf_spine_ow_I[5].z ;
 wire \tbuf_spine_ow_I[6].z ;
 wire \tbuf_spine_ow_I[7].z ;
 wire \tbuf_spine_ow_I[8].z ;
 wire \tbuf_spine_ow_I[9].z ;
 wire \zbuf_bus_iw_I[0].genblk1.l ;
 wire \zbuf_bus_iw_I[10].genblk1.l ;
 wire \zbuf_bus_iw_I[11].genblk1.l ;
 wire \zbuf_bus_iw_I[12].genblk1.l ;
 wire \zbuf_bus_iw_I[13].genblk1.l ;
 wire \zbuf_bus_iw_I[14].genblk1.l ;
 wire \zbuf_bus_iw_I[15].genblk1.l ;
 wire \zbuf_bus_iw_I[16].genblk1.l ;
 wire \zbuf_bus_iw_I[17].genblk1.l ;
 wire \zbuf_bus_iw_I[1].genblk1.l ;
 wire \zbuf_bus_iw_I[2].genblk1.l ;
 wire \zbuf_bus_iw_I[3].genblk1.l ;
 wire \zbuf_bus_iw_I[4].genblk1.l ;
 wire \zbuf_bus_iw_I[5].genblk1.l ;
 wire \zbuf_bus_iw_I[6].genblk1.l ;
 wire \zbuf_bus_iw_I[7].genblk1.l ;
 wire \zbuf_bus_iw_I[8].genblk1.l ;
 wire \zbuf_bus_iw_I[9].genblk1.l ;

 sg13g2_inv_1 _14_ (.Y(_00_),
    .A(\buf_bus_sel_I[3].z ));
 sg13g2_inv_1 _15_ (.Y(_01_),
    .A(\buf_bus_sel_I[2].z ));
 sg13g2_nand2b_1 _16_ (.Y(_02_),
    .B(\buf_bus_ena_I.z ),
    .A_N(\buf_bus_sel_I[4].z ));
 sg13g2_nor3_1 _17_ (.A(\buf_bus_sel_I[3].z ),
    .B(_01_),
    .C(_02_),
    .Y(\block[4].genblk1.grp_sel_buf_I.a ));
 sg13g2_nor2_1 _18_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .Y(_03_));
 sg13g2_and2_1 _19_ (.A(\block[4].genblk1.grp_sel_buf_I.z ),
    .B(_03_),
    .X(\block[4].l_ena_0_I.a ));
 sg13g2_nor2b_1 _20_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B_N(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .Y(_04_));
 sg13g2_and2_1 _21_ (.A(\block[4].genblk1.grp_sel_buf_I.z ),
    .B(_04_),
    .X(\block[5].l_ena_0_I.a ));
 sg13g2_nor2b_1 _22_ (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .B_N(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .Y(_05_));
 sg13g2_and2_1 _23_ (.A(\block[4].genblk1.grp_sel_buf_I.z ),
    .B(_05_),
    .X(\block[6].l_ena_0_I.a ));
 sg13g2_and2_1 _24_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .X(_06_));
 sg13g2_and2_1 _25_ (.A(\block[4].genblk1.grp_sel_buf_I.z ),
    .B(_06_),
    .X(\block[7].l_ena_0_I.a ));
 sg13g2_nor3_1 _26_ (.A(_00_),
    .B(\buf_bus_sel_I[2].z ),
    .C(_02_),
    .Y(\block[8].genblk1.grp_sel_buf_I.a ));
 sg13g2_and2_1 _27_ (.A(\block[8].genblk1.grp_sel_buf_I.z ),
    .B(_03_),
    .X(\block[8].l_ena_0_I.a ));
 sg13g2_and2_1 _28_ (.A(\block[8].genblk1.grp_sel_buf_I.z ),
    .B(_04_),
    .X(\block[9].l_ena_0_I.a ));
 sg13g2_and2_1 _29_ (.A(\block[8].genblk1.grp_sel_buf_I.z ),
    .B(_05_),
    .X(\block[10].l_ena_0_I.a ));
 sg13g2_and2_1 _30_ (.A(\block[8].genblk1.grp_sel_buf_I.z ),
    .B(_06_),
    .X(\block[11].l_ena_0_I.a ));
 sg13g2_nor2b_1 _31_ (.A(addr[1]),
    .B_N(\branch_addr_match_buf_I[1].z ),
    .Y(_07_));
 sg13g2_nor2b_1 _32_ (.A(\branch_addr_match_buf_I[2].z ),
    .B_N(addr[2]),
    .Y(_08_));
 sg13g2_xnor2_1 _33_ (.Y(_09_),
    .A(\branch_addr_match_buf_I[3].z ),
    .B(addr[3]));
 sg13g2_nand2b_1 _34_ (.Y(_10_),
    .B(addr[1]),
    .A_N(\branch_addr_match_buf_I[1].z ));
 sg13g2_nor2b_1 _35_ (.A(addr[2]),
    .B_N(\branch_addr_match_buf_I[2].z ),
    .Y(_11_));
 sg13g2_xnor2_1 _36_ (.Y(_12_),
    .A(\branch_addr_match_buf_I[0].z ),
    .B(addr[0]));
 sg13g2_nand4_1 _37_ (.B(_09_),
    .C(_10_),
    .A(\branch_ena_buf_I.z ),
    .Y(_13_),
    .D(_12_));
 sg13g2_nor4_1 _38_ (.A(_07_),
    .B(_08_),
    .C(_11_),
    .D(_13_),
    .Y(\branch_sel_buf_I.a ));
 sg13g2_nor3_1 _39_ (.A(\buf_bus_sel_I[3].z ),
    .B(\buf_bus_sel_I[2].z ),
    .C(_02_),
    .Y(\block[0].genblk1.grp_sel_buf_I.a ));
 sg13g2_and2_1 _40_ (.A(\block[0].genblk1.grp_sel_buf_I.z ),
    .B(_03_),
    .X(\block[0].l_ena_0_I.a ));
 sg13g2_and2_1 _41_ (.A(\block[0].genblk1.grp_sel_buf_I.z ),
    .B(_04_),
    .X(\block[1].l_ena_0_I.a ));
 sg13g2_and2_1 _42_ (.A(\block[0].genblk1.grp_sel_buf_I.z ),
    .B(_05_),
    .X(\block[2].l_ena_0_I.a ));
 sg13g2_and2_1 _43_ (.A(\block[0].genblk1.grp_sel_buf_I.z ),
    .B(_06_),
    .X(\block[3].l_ena_0_I.a ));
 sg13g2_antennanp \block[0].diode_I[0].cell0_I  (.A(um_ow[0]));
 sg13g2_antennanp \block[0].diode_I[10].cell0_I  (.A(um_ow[10]));
 sg13g2_antennanp \block[0].diode_I[11].cell0_I  (.A(um_ow[11]));
 sg13g2_antennanp \block[0].diode_I[12].cell0_I  (.A(um_ow[12]));
 sg13g2_antennanp \block[0].diode_I[13].cell0_I  (.A(um_ow[13]));
 sg13g2_antennanp \block[0].diode_I[14].cell0_I  (.A(um_ow[14]));
 sg13g2_antennanp \block[0].diode_I[15].cell0_I  (.A(um_ow[15]));
 sg13g2_antennanp \block[0].diode_I[16].cell0_I  (.A(um_ow[16]));
 sg13g2_antennanp \block[0].diode_I[17].cell0_I  (.A(um_ow[17]));
 sg13g2_antennanp \block[0].diode_I[18].cell0_I  (.A(um_ow[18]));
 sg13g2_antennanp \block[0].diode_I[19].cell0_I  (.A(um_ow[19]));
 sg13g2_antennanp \block[0].diode_I[1].cell0_I  (.A(um_ow[1]));
 sg13g2_antennanp \block[0].diode_I[20].cell0_I  (.A(um_ow[20]));
 sg13g2_antennanp \block[0].diode_I[21].cell0_I  (.A(um_ow[21]));
 sg13g2_antennanp \block[0].diode_I[22].cell0_I  (.A(um_ow[22]));
 sg13g2_antennanp \block[0].diode_I[23].cell0_I  (.A(um_ow[23]));
 sg13g2_antennanp \block[0].diode_I[2].cell0_I  (.A(um_ow[2]));
 sg13g2_antennanp \block[0].diode_I[3].cell0_I  (.A(um_ow[3]));
 sg13g2_antennanp \block[0].diode_I[4].cell0_I  (.A(um_ow[4]));
 sg13g2_antennanp \block[0].diode_I[5].cell0_I  (.A(um_ow[5]));
 sg13g2_antennanp \block[0].diode_I[6].cell0_I  (.A(um_ow[6]));
 sg13g2_antennanp \block[0].diode_I[7].cell0_I  (.A(um_ow[7]));
 sg13g2_antennanp \block[0].diode_I[8].cell0_I  (.A(um_ow[8]));
 sg13g2_antennanp \block[0].diode_I[9].cell0_I  (.A(um_ow[9]));
 sg13g2_buf_2 \block[0].genblk1.grp_sel_buf_I.genblk1.cell0_I  (.A(\block[0].genblk1.grp_sel_buf_I.a ),
    .X(\block[0].genblk1.grp_sel_buf_I.z ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[0].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[0]),
    .A1(um_ow[24]),
    .A2(um_ow[48]),
    .A3(um_ow[72]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[0].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[10].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[10]),
    .A1(um_ow[34]),
    .A2(um_ow[58]),
    .A3(um_ow[82]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[10].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[11].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[11]),
    .A1(um_ow[35]),
    .A2(um_ow[59]),
    .A3(um_ow[83]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[11].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[12].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[12]),
    .A1(um_ow[36]),
    .A2(um_ow[60]),
    .A3(um_ow[84]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[12].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[13].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[13]),
    .A1(um_ow[37]),
    .A2(um_ow[61]),
    .A3(um_ow[85]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[13].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[14].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[14]),
    .A1(um_ow[38]),
    .A2(um_ow[62]),
    .A3(um_ow[86]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[14].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[15].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[15]),
    .A1(um_ow[39]),
    .A2(um_ow[63]),
    .A3(um_ow[87]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[15].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[16].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[16]),
    .A1(um_ow[40]),
    .A2(um_ow[64]),
    .A3(um_ow[88]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[16].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[17].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[17]),
    .A1(um_ow[41]),
    .A2(um_ow[65]),
    .A3(um_ow[89]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[17].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[18].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[18]),
    .A1(um_ow[42]),
    .A2(um_ow[66]),
    .A3(um_ow[90]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[18].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[19].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[19]),
    .A1(um_ow[43]),
    .A2(um_ow[67]),
    .A3(um_ow[91]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[19].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[1].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[1]),
    .A1(um_ow[25]),
    .A2(um_ow[49]),
    .A3(um_ow[73]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[1].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[20].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[20]),
    .A1(um_ow[44]),
    .A2(um_ow[68]),
    .A3(um_ow[92]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[20].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[21].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[21]),
    .A1(um_ow[45]),
    .A2(um_ow[69]),
    .A3(um_ow[93]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[21].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[22].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[22]),
    .A1(um_ow[46]),
    .A2(um_ow[70]),
    .A3(um_ow[94]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[22].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[23].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[23]),
    .A1(um_ow[47]),
    .A2(um_ow[71]),
    .A3(um_ow[95]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[23].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[2].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[2]),
    .A1(um_ow[26]),
    .A2(um_ow[50]),
    .A3(um_ow[74]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[2].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[3].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[3]),
    .A1(um_ow[27]),
    .A2(um_ow[51]),
    .A3(um_ow[75]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[3].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[4].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[4]),
    .A1(um_ow[28]),
    .A2(um_ow[52]),
    .A3(um_ow[76]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[4].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[5].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[5]),
    .A1(um_ow[29]),
    .A2(um_ow[53]),
    .A3(um_ow[77]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[5].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[6].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[6]),
    .A1(um_ow[30]),
    .A2(um_ow[54]),
    .A3(um_ow[78]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[6].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[7].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[7]),
    .A1(um_ow[31]),
    .A2(um_ow[55]),
    .A3(um_ow[79]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[7].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[8].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[8]),
    .A1(um_ow[32]),
    .A2(um_ow[56]),
    .A3(um_ow[80]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[8].x ));
 sg13g2_mux4_1 \block[0].genblk1.mux4_I[9].cell0_I  (.S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[9]),
    .A1(um_ow[33]),
    .A2(um_ow[57]),
    .A3(um_ow[81]),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[9].x ));
 sg13g2_buf_2 \block[0].genblk1.mux4_sel_buf_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .X(\block[0].genblk1.mux4_sel_buf_I[0].z ));
 sg13g2_buf_2 \block[0].genblk1.mux4_sel_buf_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .X(\block[0].genblk1.mux4_sel_buf_I[1].z ));
 sg13g2_inv_8 \block[0].genblk1.tbuf_blk_ena_I.cell0_I  (.Y(\block[0].genblk1.l_tbe ),
    .A(\block[0].genblk1.grp_sel_buf_I.z ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[0].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ),
    .A(\block[0].genblk1.mux4_I[0].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[10].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ),
    .A(\block[0].genblk1.mux4_I[10].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[11].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ),
    .A(\block[0].genblk1.mux4_I[11].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[12].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ),
    .A(\block[0].genblk1.mux4_I[12].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[13].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ),
    .A(\block[0].genblk1.mux4_I[13].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[14].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ),
    .A(\block[0].genblk1.mux4_I[14].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[15].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ),
    .A(\block[0].genblk1.mux4_I[15].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[16].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ),
    .A(\block[0].genblk1.mux4_I[16].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[17].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ),
    .A(\block[0].genblk1.mux4_I[17].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[18].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ),
    .A(\block[0].genblk1.mux4_I[18].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[19].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ),
    .A(\block[0].genblk1.mux4_I[19].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[1].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ),
    .A(\block[0].genblk1.mux4_I[1].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[20].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ),
    .A(\block[0].genblk1.mux4_I[20].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[21].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ),
    .A(\block[0].genblk1.mux4_I[21].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[22].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ),
    .A(\block[0].genblk1.mux4_I[22].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[23].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ),
    .A(\block[0].genblk1.mux4_I[23].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[2].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ),
    .A(\block[0].genblk1.mux4_I[2].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[3].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ),
    .A(\block[0].genblk1.mux4_I[3].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[4].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ),
    .A(\block[0].genblk1.mux4_I[4].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[5].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ),
    .A(\block[0].genblk1.mux4_I[5].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[6].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ),
    .A(\block[0].genblk1.mux4_I[6].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[7].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ),
    .A(\block[0].genblk1.mux4_I[7].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[8].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ),
    .A(\block[0].genblk1.mux4_I[8].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[9].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ),
    .A(\block[0].genblk1.mux4_I[9].x ),
    .TE_B(\block[0].genblk1.l_tbe ));
 sg13g2_buf_8 \block[0].l_ena_0_I.genblk1.cell0_I  (.A(\block[0].l_ena_0_I.a ),
    .X(\block[0].l_ena ));
 sg13g2_tielo \block[0].tie_I.genblk1.cell0_I  (.L_LO(\block[0].tie_I.lo ));
 sg13g2_buf_2 \block[0].zbuf_ena_I.genblk1.cell0_I  (.A(\block[0].l_ena ),
    .X(\block[0].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[0].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[0].l_ena ),
    .X(\block[0].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[0].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[0].l_ena ),
    .X(\block[0].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[10].diode_I[0].cell0_I  (.A(um_ow[240]));
 sg13g2_antennanp \block[10].diode_I[10].cell0_I  (.A(um_ow[250]));
 sg13g2_antennanp \block[10].diode_I[11].cell0_I  (.A(um_ow[251]));
 sg13g2_antennanp \block[10].diode_I[12].cell0_I  (.A(um_ow[252]));
 sg13g2_antennanp \block[10].diode_I[13].cell0_I  (.A(um_ow[253]));
 sg13g2_antennanp \block[10].diode_I[14].cell0_I  (.A(um_ow[254]));
 sg13g2_antennanp \block[10].diode_I[15].cell0_I  (.A(um_ow[255]));
 sg13g2_antennanp \block[10].diode_I[16].cell0_I  (.A(um_ow[256]));
 sg13g2_antennanp \block[10].diode_I[17].cell0_I  (.A(um_ow[257]));
 sg13g2_antennanp \block[10].diode_I[18].cell0_I  (.A(um_ow[258]));
 sg13g2_antennanp \block[10].diode_I[19].cell0_I  (.A(um_ow[259]));
 sg13g2_antennanp \block[10].diode_I[1].cell0_I  (.A(um_ow[241]));
 sg13g2_antennanp \block[10].diode_I[20].cell0_I  (.A(um_ow[260]));
 sg13g2_antennanp \block[10].diode_I[21].cell0_I  (.A(um_ow[261]));
 sg13g2_antennanp \block[10].diode_I[22].cell0_I  (.A(um_ow[262]));
 sg13g2_antennanp \block[10].diode_I[23].cell0_I  (.A(um_ow[263]));
 sg13g2_antennanp \block[10].diode_I[2].cell0_I  (.A(um_ow[242]));
 sg13g2_antennanp \block[10].diode_I[3].cell0_I  (.A(um_ow[243]));
 sg13g2_antennanp \block[10].diode_I[4].cell0_I  (.A(um_ow[244]));
 sg13g2_antennanp \block[10].diode_I[5].cell0_I  (.A(um_ow[245]));
 sg13g2_antennanp \block[10].diode_I[6].cell0_I  (.A(um_ow[246]));
 sg13g2_antennanp \block[10].diode_I[7].cell0_I  (.A(um_ow[247]));
 sg13g2_antennanp \block[10].diode_I[8].cell0_I  (.A(um_ow[248]));
 sg13g2_antennanp \block[10].diode_I[9].cell0_I  (.A(um_ow[249]));
 sg13g2_buf_8 \block[10].l_ena_0_I.genblk1.cell0_I  (.A(\block[10].l_ena_0_I.a ),
    .X(\block[10].l_ena ));
 sg13g2_tielo \block[10].tie_I.genblk1.cell0_I  (.L_LO(\block[10].tie_I.lo ));
 sg13g2_buf_2 \block[10].zbuf_ena_I.genblk1.cell0_I  (.A(\block[10].l_ena ),
    .X(\block[10].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[10].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[10].l_ena ),
    .X(\block[10].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[10].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[10].l_ena ),
    .X(\block[10].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[11].diode_I[0].cell0_I  (.A(um_ow[264]));
 sg13g2_antennanp \block[11].diode_I[10].cell0_I  (.A(um_ow[274]));
 sg13g2_antennanp \block[11].diode_I[11].cell0_I  (.A(um_ow[275]));
 sg13g2_antennanp \block[11].diode_I[12].cell0_I  (.A(um_ow[276]));
 sg13g2_antennanp \block[11].diode_I[13].cell0_I  (.A(um_ow[277]));
 sg13g2_antennanp \block[11].diode_I[14].cell0_I  (.A(um_ow[278]));
 sg13g2_antennanp \block[11].diode_I[15].cell0_I  (.A(um_ow[279]));
 sg13g2_antennanp \block[11].diode_I[16].cell0_I  (.A(um_ow[280]));
 sg13g2_antennanp \block[11].diode_I[17].cell0_I  (.A(um_ow[281]));
 sg13g2_antennanp \block[11].diode_I[18].cell0_I  (.A(um_ow[282]));
 sg13g2_antennanp \block[11].diode_I[19].cell0_I  (.A(um_ow[283]));
 sg13g2_antennanp \block[11].diode_I[1].cell0_I  (.A(um_ow[265]));
 sg13g2_antennanp \block[11].diode_I[20].cell0_I  (.A(um_ow[284]));
 sg13g2_antennanp \block[11].diode_I[21].cell0_I  (.A(um_ow[285]));
 sg13g2_antennanp \block[11].diode_I[22].cell0_I  (.A(um_ow[286]));
 sg13g2_antennanp \block[11].diode_I[23].cell0_I  (.A(um_ow[287]));
 sg13g2_antennanp \block[11].diode_I[2].cell0_I  (.A(um_ow[266]));
 sg13g2_antennanp \block[11].diode_I[3].cell0_I  (.A(um_ow[267]));
 sg13g2_antennanp \block[11].diode_I[4].cell0_I  (.A(um_ow[268]));
 sg13g2_antennanp \block[11].diode_I[5].cell0_I  (.A(um_ow[269]));
 sg13g2_antennanp \block[11].diode_I[6].cell0_I  (.A(um_ow[270]));
 sg13g2_antennanp \block[11].diode_I[7].cell0_I  (.A(um_ow[271]));
 sg13g2_antennanp \block[11].diode_I[8].cell0_I  (.A(um_ow[272]));
 sg13g2_antennanp \block[11].diode_I[9].cell0_I  (.A(um_ow[273]));
 sg13g2_buf_8 \block[11].l_ena_0_I.genblk1.cell0_I  (.A(\block[11].l_ena_0_I.a ),
    .X(\block[11].l_ena ));
 sg13g2_tielo \block[11].tie_I.genblk1.cell0_I  (.L_LO(\block[11].tie_I.lo ));
 sg13g2_buf_2 \block[11].zbuf_ena_I.genblk1.cell0_I  (.A(\block[11].l_ena ),
    .X(\block[11].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[11].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[11].l_ena ),
    .X(\block[11].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[11].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[11].l_ena ),
    .X(\block[11].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[1].diode_I[0].cell0_I  (.A(um_ow[24]));
 sg13g2_antennanp \block[1].diode_I[10].cell0_I  (.A(um_ow[34]));
 sg13g2_antennanp \block[1].diode_I[11].cell0_I  (.A(um_ow[35]));
 sg13g2_antennanp \block[1].diode_I[12].cell0_I  (.A(um_ow[36]));
 sg13g2_antennanp \block[1].diode_I[13].cell0_I  (.A(um_ow[37]));
 sg13g2_antennanp \block[1].diode_I[14].cell0_I  (.A(um_ow[38]));
 sg13g2_antennanp \block[1].diode_I[15].cell0_I  (.A(um_ow[39]));
 sg13g2_antennanp \block[1].diode_I[16].cell0_I  (.A(um_ow[40]));
 sg13g2_antennanp \block[1].diode_I[17].cell0_I  (.A(um_ow[41]));
 sg13g2_antennanp \block[1].diode_I[18].cell0_I  (.A(um_ow[42]));
 sg13g2_antennanp \block[1].diode_I[19].cell0_I  (.A(um_ow[43]));
 sg13g2_antennanp \block[1].diode_I[1].cell0_I  (.A(um_ow[25]));
 sg13g2_antennanp \block[1].diode_I[20].cell0_I  (.A(um_ow[44]));
 sg13g2_antennanp \block[1].diode_I[21].cell0_I  (.A(um_ow[45]));
 sg13g2_antennanp \block[1].diode_I[22].cell0_I  (.A(um_ow[46]));
 sg13g2_antennanp \block[1].diode_I[23].cell0_I  (.A(um_ow[47]));
 sg13g2_antennanp \block[1].diode_I[2].cell0_I  (.A(um_ow[26]));
 sg13g2_antennanp \block[1].diode_I[3].cell0_I  (.A(um_ow[27]));
 sg13g2_antennanp \block[1].diode_I[4].cell0_I  (.A(um_ow[28]));
 sg13g2_antennanp \block[1].diode_I[5].cell0_I  (.A(um_ow[29]));
 sg13g2_antennanp \block[1].diode_I[6].cell0_I  (.A(um_ow[30]));
 sg13g2_antennanp \block[1].diode_I[7].cell0_I  (.A(um_ow[31]));
 sg13g2_antennanp \block[1].diode_I[8].cell0_I  (.A(um_ow[32]));
 sg13g2_antennanp \block[1].diode_I[9].cell0_I  (.A(um_ow[33]));
 sg13g2_buf_8 \block[1].l_ena_0_I.genblk1.cell0_I  (.A(\block[1].l_ena_0_I.a ),
    .X(\block[1].l_ena ));
 sg13g2_tielo \block[1].tie_I.genblk1.cell0_I  (.L_LO(\block[1].tie_I.lo ));
 sg13g2_buf_2 \block[1].zbuf_ena_I.genblk1.cell0_I  (.A(\block[1].l_ena ),
    .X(\block[1].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[1].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[1].l_ena ),
    .X(\block[1].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[1].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[1].l_ena ),
    .X(\block[1].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[2].diode_I[0].cell0_I  (.A(um_ow[48]));
 sg13g2_antennanp \block[2].diode_I[10].cell0_I  (.A(um_ow[58]));
 sg13g2_antennanp \block[2].diode_I[11].cell0_I  (.A(um_ow[59]));
 sg13g2_antennanp \block[2].diode_I[12].cell0_I  (.A(um_ow[60]));
 sg13g2_antennanp \block[2].diode_I[13].cell0_I  (.A(um_ow[61]));
 sg13g2_antennanp \block[2].diode_I[14].cell0_I  (.A(um_ow[62]));
 sg13g2_antennanp \block[2].diode_I[15].cell0_I  (.A(um_ow[63]));
 sg13g2_antennanp \block[2].diode_I[16].cell0_I  (.A(um_ow[64]));
 sg13g2_antennanp \block[2].diode_I[17].cell0_I  (.A(um_ow[65]));
 sg13g2_antennanp \block[2].diode_I[18].cell0_I  (.A(um_ow[66]));
 sg13g2_antennanp \block[2].diode_I[19].cell0_I  (.A(um_ow[67]));
 sg13g2_antennanp \block[2].diode_I[1].cell0_I  (.A(um_ow[49]));
 sg13g2_antennanp \block[2].diode_I[20].cell0_I  (.A(um_ow[68]));
 sg13g2_antennanp \block[2].diode_I[21].cell0_I  (.A(um_ow[69]));
 sg13g2_antennanp \block[2].diode_I[22].cell0_I  (.A(um_ow[70]));
 sg13g2_antennanp \block[2].diode_I[23].cell0_I  (.A(um_ow[71]));
 sg13g2_antennanp \block[2].diode_I[2].cell0_I  (.A(um_ow[50]));
 sg13g2_antennanp \block[2].diode_I[3].cell0_I  (.A(um_ow[51]));
 sg13g2_antennanp \block[2].diode_I[4].cell0_I  (.A(um_ow[52]));
 sg13g2_antennanp \block[2].diode_I[5].cell0_I  (.A(um_ow[53]));
 sg13g2_antennanp \block[2].diode_I[6].cell0_I  (.A(um_ow[54]));
 sg13g2_antennanp \block[2].diode_I[7].cell0_I  (.A(um_ow[55]));
 sg13g2_antennanp \block[2].diode_I[8].cell0_I  (.A(um_ow[56]));
 sg13g2_antennanp \block[2].diode_I[9].cell0_I  (.A(um_ow[57]));
 sg13g2_buf_8 \block[2].l_ena_0_I.genblk1.cell0_I  (.A(\block[2].l_ena_0_I.a ),
    .X(\block[2].l_ena ));
 sg13g2_tielo \block[2].tie_I.genblk1.cell0_I  (.L_LO(\block[2].tie_I.lo ));
 sg13g2_buf_2 \block[2].zbuf_ena_I.genblk1.cell0_I  (.A(\block[2].l_ena ),
    .X(\block[2].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[2].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[2].l_ena ),
    .X(\block[2].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[2].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[2].l_ena ),
    .X(\block[2].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[3].diode_I[0].cell0_I  (.A(um_ow[72]));
 sg13g2_antennanp \block[3].diode_I[10].cell0_I  (.A(um_ow[82]));
 sg13g2_antennanp \block[3].diode_I[11].cell0_I  (.A(um_ow[83]));
 sg13g2_antennanp \block[3].diode_I[12].cell0_I  (.A(um_ow[84]));
 sg13g2_antennanp \block[3].diode_I[13].cell0_I  (.A(um_ow[85]));
 sg13g2_antennanp \block[3].diode_I[14].cell0_I  (.A(um_ow[86]));
 sg13g2_antennanp \block[3].diode_I[15].cell0_I  (.A(um_ow[87]));
 sg13g2_antennanp \block[3].diode_I[16].cell0_I  (.A(um_ow[88]));
 sg13g2_antennanp \block[3].diode_I[17].cell0_I  (.A(um_ow[89]));
 sg13g2_antennanp \block[3].diode_I[18].cell0_I  (.A(um_ow[90]));
 sg13g2_antennanp \block[3].diode_I[19].cell0_I  (.A(um_ow[91]));
 sg13g2_antennanp \block[3].diode_I[1].cell0_I  (.A(um_ow[73]));
 sg13g2_antennanp \block[3].diode_I[20].cell0_I  (.A(um_ow[92]));
 sg13g2_antennanp \block[3].diode_I[21].cell0_I  (.A(um_ow[93]));
 sg13g2_antennanp \block[3].diode_I[22].cell0_I  (.A(um_ow[94]));
 sg13g2_antennanp \block[3].diode_I[23].cell0_I  (.A(um_ow[95]));
 sg13g2_antennanp \block[3].diode_I[2].cell0_I  (.A(um_ow[74]));
 sg13g2_antennanp \block[3].diode_I[3].cell0_I  (.A(um_ow[75]));
 sg13g2_antennanp \block[3].diode_I[4].cell0_I  (.A(um_ow[76]));
 sg13g2_antennanp \block[3].diode_I[5].cell0_I  (.A(um_ow[77]));
 sg13g2_antennanp \block[3].diode_I[6].cell0_I  (.A(um_ow[78]));
 sg13g2_antennanp \block[3].diode_I[7].cell0_I  (.A(um_ow[79]));
 sg13g2_antennanp \block[3].diode_I[8].cell0_I  (.A(um_ow[80]));
 sg13g2_antennanp \block[3].diode_I[9].cell0_I  (.A(um_ow[81]));
 sg13g2_buf_8 \block[3].l_ena_0_I.genblk1.cell0_I  (.A(\block[3].l_ena_0_I.a ),
    .X(\block[3].l_ena ));
 sg13g2_tielo \block[3].tie_I.genblk1.cell0_I  (.L_LO(\block[3].tie_I.lo ));
 sg13g2_buf_2 \block[3].zbuf_ena_I.genblk1.cell0_I  (.A(\block[3].l_ena ),
    .X(\block[3].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[3].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[3].l_ena ),
    .X(\block[3].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[3].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[3].l_ena ),
    .X(\block[3].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[4].diode_I[0].cell0_I  (.A(um_ow[96]));
 sg13g2_antennanp \block[4].diode_I[10].cell0_I  (.A(um_ow[106]));
 sg13g2_antennanp \block[4].diode_I[11].cell0_I  (.A(um_ow[107]));
 sg13g2_antennanp \block[4].diode_I[12].cell0_I  (.A(um_ow[108]));
 sg13g2_antennanp \block[4].diode_I[13].cell0_I  (.A(um_ow[109]));
 sg13g2_antennanp \block[4].diode_I[14].cell0_I  (.A(um_ow[110]));
 sg13g2_antennanp \block[4].diode_I[15].cell0_I  (.A(um_ow[111]));
 sg13g2_antennanp \block[4].diode_I[16].cell0_I  (.A(um_ow[112]));
 sg13g2_antennanp \block[4].diode_I[17].cell0_I  (.A(um_ow[113]));
 sg13g2_antennanp \block[4].diode_I[18].cell0_I  (.A(um_ow[114]));
 sg13g2_antennanp \block[4].diode_I[19].cell0_I  (.A(um_ow[115]));
 sg13g2_antennanp \block[4].diode_I[1].cell0_I  (.A(um_ow[97]));
 sg13g2_antennanp \block[4].diode_I[20].cell0_I  (.A(um_ow[116]));
 sg13g2_antennanp \block[4].diode_I[21].cell0_I  (.A(um_ow[117]));
 sg13g2_antennanp \block[4].diode_I[22].cell0_I  (.A(um_ow[118]));
 sg13g2_antennanp \block[4].diode_I[23].cell0_I  (.A(um_ow[119]));
 sg13g2_antennanp \block[4].diode_I[2].cell0_I  (.A(um_ow[98]));
 sg13g2_antennanp \block[4].diode_I[3].cell0_I  (.A(um_ow[99]));
 sg13g2_antennanp \block[4].diode_I[4].cell0_I  (.A(um_ow[100]));
 sg13g2_antennanp \block[4].diode_I[5].cell0_I  (.A(um_ow[101]));
 sg13g2_antennanp \block[4].diode_I[6].cell0_I  (.A(um_ow[102]));
 sg13g2_antennanp \block[4].diode_I[7].cell0_I  (.A(um_ow[103]));
 sg13g2_antennanp \block[4].diode_I[8].cell0_I  (.A(um_ow[104]));
 sg13g2_antennanp \block[4].diode_I[9].cell0_I  (.A(um_ow[105]));
 sg13g2_buf_2 \block[4].genblk1.grp_sel_buf_I.genblk1.cell0_I  (.A(\block[4].genblk1.grp_sel_buf_I.a ),
    .X(\block[4].genblk1.grp_sel_buf_I.z ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[0].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[96]),
    .A1(um_ow[120]),
    .A2(um_ow[144]),
    .A3(um_ow[168]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[0].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[10].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[106]),
    .A1(um_ow[130]),
    .A2(um_ow[154]),
    .A3(um_ow[178]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[10].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[11].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[107]),
    .A1(um_ow[131]),
    .A2(um_ow[155]),
    .A3(um_ow[179]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[11].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[12].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[108]),
    .A1(um_ow[132]),
    .A2(um_ow[156]),
    .A3(um_ow[180]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[12].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[13].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[109]),
    .A1(um_ow[133]),
    .A2(um_ow[157]),
    .A3(um_ow[181]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[13].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[14].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[110]),
    .A1(um_ow[134]),
    .A2(um_ow[158]),
    .A3(um_ow[182]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[14].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[15].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[111]),
    .A1(um_ow[135]),
    .A2(um_ow[159]),
    .A3(um_ow[183]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[15].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[16].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[112]),
    .A1(um_ow[136]),
    .A2(um_ow[160]),
    .A3(um_ow[184]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[16].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[17].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[113]),
    .A1(um_ow[137]),
    .A2(um_ow[161]),
    .A3(um_ow[185]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[17].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[18].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[114]),
    .A1(um_ow[138]),
    .A2(um_ow[162]),
    .A3(um_ow[186]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[18].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[19].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[115]),
    .A1(um_ow[139]),
    .A2(um_ow[163]),
    .A3(um_ow[187]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[19].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[1].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[97]),
    .A1(um_ow[121]),
    .A2(um_ow[145]),
    .A3(um_ow[169]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[1].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[20].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[116]),
    .A1(um_ow[140]),
    .A2(um_ow[164]),
    .A3(um_ow[188]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[20].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[21].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[117]),
    .A1(um_ow[141]),
    .A2(um_ow[165]),
    .A3(um_ow[189]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[21].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[22].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[118]),
    .A1(um_ow[142]),
    .A2(um_ow[166]),
    .A3(um_ow[190]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[22].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[23].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[119]),
    .A1(um_ow[143]),
    .A2(um_ow[167]),
    .A3(um_ow[191]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[23].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[2].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[98]),
    .A1(um_ow[122]),
    .A2(um_ow[146]),
    .A3(um_ow[170]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[2].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[3].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[99]),
    .A1(um_ow[123]),
    .A2(um_ow[147]),
    .A3(um_ow[171]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[3].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[4].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[100]),
    .A1(um_ow[124]),
    .A2(um_ow[148]),
    .A3(um_ow[172]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[4].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[5].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[101]),
    .A1(um_ow[125]),
    .A2(um_ow[149]),
    .A3(um_ow[173]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[5].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[6].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[102]),
    .A1(um_ow[126]),
    .A2(um_ow[150]),
    .A3(um_ow[174]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[6].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[7].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[103]),
    .A1(um_ow[127]),
    .A2(um_ow[151]),
    .A3(um_ow[175]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[7].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[8].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[104]),
    .A1(um_ow[128]),
    .A2(um_ow[152]),
    .A3(um_ow[176]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[8].x ));
 sg13g2_mux4_1 \block[4].genblk1.mux4_I[9].cell0_I  (.S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[105]),
    .A1(um_ow[129]),
    .A2(um_ow[153]),
    .A3(um_ow[177]),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[9].x ));
 sg13g2_buf_2 \block[4].genblk1.mux4_sel_buf_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .X(\block[4].genblk1.mux4_sel_buf_I[0].z ));
 sg13g2_buf_2 \block[4].genblk1.mux4_sel_buf_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .X(\block[4].genblk1.mux4_sel_buf_I[1].z ));
 sg13g2_inv_8 \block[4].genblk1.tbuf_blk_ena_I.cell0_I  (.Y(\block[4].genblk1.l_tbe ),
    .A(\block[4].genblk1.grp_sel_buf_I.z ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[0].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ),
    .A(\block[4].genblk1.mux4_I[0].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[10].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ),
    .A(\block[4].genblk1.mux4_I[10].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[11].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ),
    .A(\block[4].genblk1.mux4_I[11].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[12].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ),
    .A(\block[4].genblk1.mux4_I[12].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[13].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ),
    .A(\block[4].genblk1.mux4_I[13].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[14].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ),
    .A(\block[4].genblk1.mux4_I[14].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[15].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ),
    .A(\block[4].genblk1.mux4_I[15].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[16].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ),
    .A(\block[4].genblk1.mux4_I[16].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[17].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ),
    .A(\block[4].genblk1.mux4_I[17].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[18].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ),
    .A(\block[4].genblk1.mux4_I[18].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[19].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ),
    .A(\block[4].genblk1.mux4_I[19].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[1].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ),
    .A(\block[4].genblk1.mux4_I[1].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[20].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ),
    .A(\block[4].genblk1.mux4_I[20].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[21].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ),
    .A(\block[4].genblk1.mux4_I[21].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[22].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ),
    .A(\block[4].genblk1.mux4_I[22].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[23].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ),
    .A(\block[4].genblk1.mux4_I[23].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[2].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ),
    .A(\block[4].genblk1.mux4_I[2].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[3].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ),
    .A(\block[4].genblk1.mux4_I[3].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[4].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ),
    .A(\block[4].genblk1.mux4_I[4].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[5].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ),
    .A(\block[4].genblk1.mux4_I[5].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[6].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ),
    .A(\block[4].genblk1.mux4_I[6].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[7].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ),
    .A(\block[4].genblk1.mux4_I[7].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[8].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ),
    .A(\block[4].genblk1.mux4_I[8].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[9].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ),
    .A(\block[4].genblk1.mux4_I[9].x ),
    .TE_B(\block[4].genblk1.l_tbe ));
 sg13g2_buf_8 \block[4].l_ena_0_I.genblk1.cell0_I  (.A(\block[4].l_ena_0_I.a ),
    .X(\block[4].l_ena ));
 sg13g2_tielo \block[4].tie_I.genblk1.cell0_I  (.L_LO(\block[4].tie_I.lo ));
 sg13g2_buf_2 \block[4].zbuf_ena_I.genblk1.cell0_I  (.A(\block[4].l_ena ),
    .X(\block[4].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[4].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[4].l_ena ),
    .X(\block[4].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[4].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[4].l_ena ),
    .X(\block[4].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[5].diode_I[0].cell0_I  (.A(um_ow[120]));
 sg13g2_antennanp \block[5].diode_I[10].cell0_I  (.A(um_ow[130]));
 sg13g2_antennanp \block[5].diode_I[11].cell0_I  (.A(um_ow[131]));
 sg13g2_antennanp \block[5].diode_I[12].cell0_I  (.A(um_ow[132]));
 sg13g2_antennanp \block[5].diode_I[13].cell0_I  (.A(um_ow[133]));
 sg13g2_antennanp \block[5].diode_I[14].cell0_I  (.A(um_ow[134]));
 sg13g2_antennanp \block[5].diode_I[15].cell0_I  (.A(um_ow[135]));
 sg13g2_antennanp \block[5].diode_I[16].cell0_I  (.A(um_ow[136]));
 sg13g2_antennanp \block[5].diode_I[17].cell0_I  (.A(um_ow[137]));
 sg13g2_antennanp \block[5].diode_I[18].cell0_I  (.A(um_ow[138]));
 sg13g2_antennanp \block[5].diode_I[19].cell0_I  (.A(um_ow[139]));
 sg13g2_antennanp \block[5].diode_I[1].cell0_I  (.A(um_ow[121]));
 sg13g2_antennanp \block[5].diode_I[20].cell0_I  (.A(um_ow[140]));
 sg13g2_antennanp \block[5].diode_I[21].cell0_I  (.A(um_ow[141]));
 sg13g2_antennanp \block[5].diode_I[22].cell0_I  (.A(um_ow[142]));
 sg13g2_antennanp \block[5].diode_I[23].cell0_I  (.A(um_ow[143]));
 sg13g2_antennanp \block[5].diode_I[2].cell0_I  (.A(um_ow[122]));
 sg13g2_antennanp \block[5].diode_I[3].cell0_I  (.A(um_ow[123]));
 sg13g2_antennanp \block[5].diode_I[4].cell0_I  (.A(um_ow[124]));
 sg13g2_antennanp \block[5].diode_I[5].cell0_I  (.A(um_ow[125]));
 sg13g2_antennanp \block[5].diode_I[6].cell0_I  (.A(um_ow[126]));
 sg13g2_antennanp \block[5].diode_I[7].cell0_I  (.A(um_ow[127]));
 sg13g2_antennanp \block[5].diode_I[8].cell0_I  (.A(um_ow[128]));
 sg13g2_antennanp \block[5].diode_I[9].cell0_I  (.A(um_ow[129]));
 sg13g2_buf_8 \block[5].l_ena_0_I.genblk1.cell0_I  (.A(\block[5].l_ena_0_I.a ),
    .X(\block[5].l_ena ));
 sg13g2_tielo \block[5].tie_I.genblk1.cell0_I  (.L_LO(\block[5].tie_I.lo ));
 sg13g2_buf_2 \block[5].zbuf_ena_I.genblk1.cell0_I  (.A(\block[5].l_ena ),
    .X(\block[5].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[5].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[5].l_ena ),
    .X(\block[5].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[5].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[5].l_ena ),
    .X(\block[5].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[6].diode_I[0].cell0_I  (.A(um_ow[144]));
 sg13g2_antennanp \block[6].diode_I[10].cell0_I  (.A(um_ow[154]));
 sg13g2_antennanp \block[6].diode_I[11].cell0_I  (.A(um_ow[155]));
 sg13g2_antennanp \block[6].diode_I[12].cell0_I  (.A(um_ow[156]));
 sg13g2_antennanp \block[6].diode_I[13].cell0_I  (.A(um_ow[157]));
 sg13g2_antennanp \block[6].diode_I[14].cell0_I  (.A(um_ow[158]));
 sg13g2_antennanp \block[6].diode_I[15].cell0_I  (.A(um_ow[159]));
 sg13g2_antennanp \block[6].diode_I[16].cell0_I  (.A(um_ow[160]));
 sg13g2_antennanp \block[6].diode_I[17].cell0_I  (.A(um_ow[161]));
 sg13g2_antennanp \block[6].diode_I[18].cell0_I  (.A(um_ow[162]));
 sg13g2_antennanp \block[6].diode_I[19].cell0_I  (.A(um_ow[163]));
 sg13g2_antennanp \block[6].diode_I[1].cell0_I  (.A(um_ow[145]));
 sg13g2_antennanp \block[6].diode_I[20].cell0_I  (.A(um_ow[164]));
 sg13g2_antennanp \block[6].diode_I[21].cell0_I  (.A(um_ow[165]));
 sg13g2_antennanp \block[6].diode_I[22].cell0_I  (.A(um_ow[166]));
 sg13g2_antennanp \block[6].diode_I[23].cell0_I  (.A(um_ow[167]));
 sg13g2_antennanp \block[6].diode_I[2].cell0_I  (.A(um_ow[146]));
 sg13g2_antennanp \block[6].diode_I[3].cell0_I  (.A(um_ow[147]));
 sg13g2_antennanp \block[6].diode_I[4].cell0_I  (.A(um_ow[148]));
 sg13g2_antennanp \block[6].diode_I[5].cell0_I  (.A(um_ow[149]));
 sg13g2_antennanp \block[6].diode_I[6].cell0_I  (.A(um_ow[150]));
 sg13g2_antennanp \block[6].diode_I[7].cell0_I  (.A(um_ow[151]));
 sg13g2_antennanp \block[6].diode_I[8].cell0_I  (.A(um_ow[152]));
 sg13g2_antennanp \block[6].diode_I[9].cell0_I  (.A(um_ow[153]));
 sg13g2_buf_8 \block[6].l_ena_0_I.genblk1.cell0_I  (.A(\block[6].l_ena_0_I.a ),
    .X(\block[6].l_ena ));
 sg13g2_tielo \block[6].tie_I.genblk1.cell0_I  (.L_LO(\block[6].tie_I.lo ));
 sg13g2_buf_2 \block[6].zbuf_ena_I.genblk1.cell0_I  (.A(\block[6].l_ena ),
    .X(\block[6].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[6].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[6].l_ena ),
    .X(\block[6].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[6].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[6].l_ena ),
    .X(\block[6].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[7].diode_I[0].cell0_I  (.A(um_ow[168]));
 sg13g2_antennanp \block[7].diode_I[10].cell0_I  (.A(um_ow[178]));
 sg13g2_antennanp \block[7].diode_I[11].cell0_I  (.A(um_ow[179]));
 sg13g2_antennanp \block[7].diode_I[12].cell0_I  (.A(um_ow[180]));
 sg13g2_antennanp \block[7].diode_I[13].cell0_I  (.A(um_ow[181]));
 sg13g2_antennanp \block[7].diode_I[14].cell0_I  (.A(um_ow[182]));
 sg13g2_antennanp \block[7].diode_I[15].cell0_I  (.A(um_ow[183]));
 sg13g2_antennanp \block[7].diode_I[16].cell0_I  (.A(um_ow[184]));
 sg13g2_antennanp \block[7].diode_I[17].cell0_I  (.A(um_ow[185]));
 sg13g2_antennanp \block[7].diode_I[18].cell0_I  (.A(um_ow[186]));
 sg13g2_antennanp \block[7].diode_I[19].cell0_I  (.A(um_ow[187]));
 sg13g2_antennanp \block[7].diode_I[1].cell0_I  (.A(um_ow[169]));
 sg13g2_antennanp \block[7].diode_I[20].cell0_I  (.A(um_ow[188]));
 sg13g2_antennanp \block[7].diode_I[21].cell0_I  (.A(um_ow[189]));
 sg13g2_antennanp \block[7].diode_I[22].cell0_I  (.A(um_ow[190]));
 sg13g2_antennanp \block[7].diode_I[23].cell0_I  (.A(um_ow[191]));
 sg13g2_antennanp \block[7].diode_I[2].cell0_I  (.A(um_ow[170]));
 sg13g2_antennanp \block[7].diode_I[3].cell0_I  (.A(um_ow[171]));
 sg13g2_antennanp \block[7].diode_I[4].cell0_I  (.A(um_ow[172]));
 sg13g2_antennanp \block[7].diode_I[5].cell0_I  (.A(um_ow[173]));
 sg13g2_antennanp \block[7].diode_I[6].cell0_I  (.A(um_ow[174]));
 sg13g2_antennanp \block[7].diode_I[7].cell0_I  (.A(um_ow[175]));
 sg13g2_antennanp \block[7].diode_I[8].cell0_I  (.A(um_ow[176]));
 sg13g2_antennanp \block[7].diode_I[9].cell0_I  (.A(um_ow[177]));
 sg13g2_buf_8 \block[7].l_ena_0_I.genblk1.cell0_I  (.A(\block[7].l_ena_0_I.a ),
    .X(\block[7].l_ena ));
 sg13g2_tielo \block[7].tie_I.genblk1.cell0_I  (.L_LO(\block[7].tie_I.lo ));
 sg13g2_buf_2 \block[7].zbuf_ena_I.genblk1.cell0_I  (.A(\block[7].l_ena ),
    .X(\block[7].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[7].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[7].l_ena ),
    .X(\block[7].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[7].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[7].l_ena ),
    .X(\block[7].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[8].diode_I[0].cell0_I  (.A(um_ow[192]));
 sg13g2_antennanp \block[8].diode_I[10].cell0_I  (.A(um_ow[202]));
 sg13g2_antennanp \block[8].diode_I[11].cell0_I  (.A(um_ow[203]));
 sg13g2_antennanp \block[8].diode_I[12].cell0_I  (.A(um_ow[204]));
 sg13g2_antennanp \block[8].diode_I[13].cell0_I  (.A(um_ow[205]));
 sg13g2_antennanp \block[8].diode_I[14].cell0_I  (.A(um_ow[206]));
 sg13g2_antennanp \block[8].diode_I[15].cell0_I  (.A(um_ow[207]));
 sg13g2_antennanp \block[8].diode_I[16].cell0_I  (.A(um_ow[208]));
 sg13g2_antennanp \block[8].diode_I[17].cell0_I  (.A(um_ow[209]));
 sg13g2_antennanp \block[8].diode_I[18].cell0_I  (.A(um_ow[210]));
 sg13g2_antennanp \block[8].diode_I[19].cell0_I  (.A(um_ow[211]));
 sg13g2_antennanp \block[8].diode_I[1].cell0_I  (.A(um_ow[193]));
 sg13g2_antennanp \block[8].diode_I[20].cell0_I  (.A(um_ow[212]));
 sg13g2_antennanp \block[8].diode_I[21].cell0_I  (.A(um_ow[213]));
 sg13g2_antennanp \block[8].diode_I[22].cell0_I  (.A(um_ow[214]));
 sg13g2_antennanp \block[8].diode_I[23].cell0_I  (.A(um_ow[215]));
 sg13g2_antennanp \block[8].diode_I[2].cell0_I  (.A(um_ow[194]));
 sg13g2_antennanp \block[8].diode_I[3].cell0_I  (.A(um_ow[195]));
 sg13g2_antennanp \block[8].diode_I[4].cell0_I  (.A(um_ow[196]));
 sg13g2_antennanp \block[8].diode_I[5].cell0_I  (.A(um_ow[197]));
 sg13g2_antennanp \block[8].diode_I[6].cell0_I  (.A(um_ow[198]));
 sg13g2_antennanp \block[8].diode_I[7].cell0_I  (.A(um_ow[199]));
 sg13g2_antennanp \block[8].diode_I[8].cell0_I  (.A(um_ow[200]));
 sg13g2_antennanp \block[8].diode_I[9].cell0_I  (.A(um_ow[201]));
 sg13g2_buf_2 \block[8].genblk1.grp_sel_buf_I.genblk1.cell0_I  (.A(\block[8].genblk1.grp_sel_buf_I.a ),
    .X(\block[8].genblk1.grp_sel_buf_I.z ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[0].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[192]),
    .A1(um_ow[216]),
    .A2(um_ow[240]),
    .A3(um_ow[264]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[0].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[10].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[202]),
    .A1(um_ow[226]),
    .A2(um_ow[250]),
    .A3(um_ow[274]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[10].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[11].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[203]),
    .A1(um_ow[227]),
    .A2(um_ow[251]),
    .A3(um_ow[275]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[11].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[12].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[204]),
    .A1(um_ow[228]),
    .A2(um_ow[252]),
    .A3(um_ow[276]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[12].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[13].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[205]),
    .A1(um_ow[229]),
    .A2(um_ow[253]),
    .A3(um_ow[277]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[13].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[14].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[206]),
    .A1(um_ow[230]),
    .A2(um_ow[254]),
    .A3(um_ow[278]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[14].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[15].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[207]),
    .A1(um_ow[231]),
    .A2(um_ow[255]),
    .A3(um_ow[279]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[15].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[16].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[208]),
    .A1(um_ow[232]),
    .A2(um_ow[256]),
    .A3(um_ow[280]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[16].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[17].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[209]),
    .A1(um_ow[233]),
    .A2(um_ow[257]),
    .A3(um_ow[281]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[17].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[18].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[210]),
    .A1(um_ow[234]),
    .A2(um_ow[258]),
    .A3(um_ow[282]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[18].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[19].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[211]),
    .A1(um_ow[235]),
    .A2(um_ow[259]),
    .A3(um_ow[283]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[19].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[1].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[193]),
    .A1(um_ow[217]),
    .A2(um_ow[241]),
    .A3(um_ow[265]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[1].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[20].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[212]),
    .A1(um_ow[236]),
    .A2(um_ow[260]),
    .A3(um_ow[284]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[20].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[21].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[213]),
    .A1(um_ow[237]),
    .A2(um_ow[261]),
    .A3(um_ow[285]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[21].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[22].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[214]),
    .A1(um_ow[238]),
    .A2(um_ow[262]),
    .A3(um_ow[286]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[22].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[23].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[215]),
    .A1(um_ow[239]),
    .A2(um_ow[263]),
    .A3(um_ow[287]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[23].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[2].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[194]),
    .A1(um_ow[218]),
    .A2(um_ow[242]),
    .A3(um_ow[266]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[2].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[3].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[195]),
    .A1(um_ow[219]),
    .A2(um_ow[243]),
    .A3(um_ow[267]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[3].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[4].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[196]),
    .A1(um_ow[220]),
    .A2(um_ow[244]),
    .A3(um_ow[268]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[4].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[5].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[197]),
    .A1(um_ow[221]),
    .A2(um_ow[245]),
    .A3(um_ow[269]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[5].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[6].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[198]),
    .A1(um_ow[222]),
    .A2(um_ow[246]),
    .A3(um_ow[270]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[6].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[7].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[199]),
    .A1(um_ow[223]),
    .A2(um_ow[247]),
    .A3(um_ow[271]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[7].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[8].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[200]),
    .A1(um_ow[224]),
    .A2(um_ow[248]),
    .A3(um_ow[272]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[8].x ));
 sg13g2_mux4_1 \block[8].genblk1.mux4_I[9].cell0_I  (.S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .A0(um_ow[201]),
    .A1(um_ow[225]),
    .A2(um_ow[249]),
    .A3(um_ow[273]),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[9].x ));
 sg13g2_buf_2 \block[8].genblk1.mux4_sel_buf_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .X(\block[8].genblk1.mux4_sel_buf_I[0].z ));
 sg13g2_buf_2 \block[8].genblk1.mux4_sel_buf_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .X(\block[8].genblk1.mux4_sel_buf_I[1].z ));
 sg13g2_inv_8 \block[8].genblk1.tbuf_blk_ena_I.cell0_I  (.Y(\block[8].genblk1.l_tbe ),
    .A(\block[8].genblk1.grp_sel_buf_I.z ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[0].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ),
    .A(\block[8].genblk1.mux4_I[0].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[10].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ),
    .A(\block[8].genblk1.mux4_I[10].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[11].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ),
    .A(\block[8].genblk1.mux4_I[11].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[12].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ),
    .A(\block[8].genblk1.mux4_I[12].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[13].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ),
    .A(\block[8].genblk1.mux4_I[13].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[14].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ),
    .A(\block[8].genblk1.mux4_I[14].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[15].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ),
    .A(\block[8].genblk1.mux4_I[15].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[16].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ),
    .A(\block[8].genblk1.mux4_I[16].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[17].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ),
    .A(\block[8].genblk1.mux4_I[17].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[18].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ),
    .A(\block[8].genblk1.mux4_I[18].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[19].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ),
    .A(\block[8].genblk1.mux4_I[19].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[1].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ),
    .A(\block[8].genblk1.mux4_I[1].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[20].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ),
    .A(\block[8].genblk1.mux4_I[20].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[21].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ),
    .A(\block[8].genblk1.mux4_I[21].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[22].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ),
    .A(\block[8].genblk1.mux4_I[22].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[23].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ),
    .A(\block[8].genblk1.mux4_I[23].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[2].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ),
    .A(\block[8].genblk1.mux4_I[2].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[3].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ),
    .A(\block[8].genblk1.mux4_I[3].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[4].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ),
    .A(\block[8].genblk1.mux4_I[4].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[5].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ),
    .A(\block[8].genblk1.mux4_I[5].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[6].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ),
    .A(\block[8].genblk1.mux4_I[6].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[7].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ),
    .A(\block[8].genblk1.mux4_I[7].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[8].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ),
    .A(\block[8].genblk1.mux4_I[8].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[9].genblk1.cell0_I  (.Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ),
    .A(\block[8].genblk1.mux4_I[9].x ),
    .TE_B(\block[8].genblk1.l_tbe ));
 sg13g2_buf_8 \block[8].l_ena_0_I.genblk1.cell0_I  (.A(\block[8].l_ena_0_I.a ),
    .X(\block[8].l_ena ));
 sg13g2_tielo \block[8].tie_I.genblk1.cell0_I  (.L_LO(\block[8].tie_I.lo ));
 sg13g2_buf_2 \block[8].zbuf_ena_I.genblk1.cell0_I  (.A(\block[8].l_ena ),
    .X(\block[8].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[8].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[8].l_ena ),
    .X(\block[8].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[8].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[8].l_ena ),
    .X(\block[8].zbuf_pg_ena_I.z ));
 sg13g2_antennanp \block[9].diode_I[0].cell0_I  (.A(um_ow[216]));
 sg13g2_antennanp \block[9].diode_I[10].cell0_I  (.A(um_ow[226]));
 sg13g2_antennanp \block[9].diode_I[11].cell0_I  (.A(um_ow[227]));
 sg13g2_antennanp \block[9].diode_I[12].cell0_I  (.A(um_ow[228]));
 sg13g2_antennanp \block[9].diode_I[13].cell0_I  (.A(um_ow[229]));
 sg13g2_antennanp \block[9].diode_I[14].cell0_I  (.A(um_ow[230]));
 sg13g2_antennanp \block[9].diode_I[15].cell0_I  (.A(um_ow[231]));
 sg13g2_antennanp \block[9].diode_I[16].cell0_I  (.A(um_ow[232]));
 sg13g2_antennanp \block[9].diode_I[17].cell0_I  (.A(um_ow[233]));
 sg13g2_antennanp \block[9].diode_I[18].cell0_I  (.A(um_ow[234]));
 sg13g2_antennanp \block[9].diode_I[19].cell0_I  (.A(um_ow[235]));
 sg13g2_antennanp \block[9].diode_I[1].cell0_I  (.A(um_ow[217]));
 sg13g2_antennanp \block[9].diode_I[20].cell0_I  (.A(um_ow[236]));
 sg13g2_antennanp \block[9].diode_I[21].cell0_I  (.A(um_ow[237]));
 sg13g2_antennanp \block[9].diode_I[22].cell0_I  (.A(um_ow[238]));
 sg13g2_antennanp \block[9].diode_I[23].cell0_I  (.A(um_ow[239]));
 sg13g2_antennanp \block[9].diode_I[2].cell0_I  (.A(um_ow[218]));
 sg13g2_antennanp \block[9].diode_I[3].cell0_I  (.A(um_ow[219]));
 sg13g2_antennanp \block[9].diode_I[4].cell0_I  (.A(um_ow[220]));
 sg13g2_antennanp \block[9].diode_I[5].cell0_I  (.A(um_ow[221]));
 sg13g2_antennanp \block[9].diode_I[6].cell0_I  (.A(um_ow[222]));
 sg13g2_antennanp \block[9].diode_I[7].cell0_I  (.A(um_ow[223]));
 sg13g2_antennanp \block[9].diode_I[8].cell0_I  (.A(um_ow[224]));
 sg13g2_antennanp \block[9].diode_I[9].cell0_I  (.A(um_ow[225]));
 sg13g2_buf_8 \block[9].l_ena_0_I.genblk1.cell0_I  (.A(\block[9].l_ena_0_I.a ),
    .X(\block[9].l_ena ));
 sg13g2_tielo \block[9].tie_I.genblk1.cell0_I  (.L_LO(\block[9].tie_I.lo ));
 sg13g2_buf_2 \block[9].zbuf_ena_I.genblk1.cell0_I  (.A(\block[9].l_ena ),
    .X(\block[9].zbuf_ena_I.z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[0].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[0].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[10].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[10].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[11].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[11].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[12].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[12].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[13].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[13].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[14].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[14].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[15].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[15].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[16].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[16].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[17].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[17].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[1].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[1].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[2].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[2].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[3].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[3].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[4].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[4].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[5].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[5].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[6].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[6].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[7].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[7].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[8].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[8].z ));
 sg13g2_and2_2 \block[9].zbuf_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_iw_I[9].a ),
    .B(\block[9].l_ena ),
    .X(\block[9].zbuf_iw_I[9].z ));
 sg13g2_buf_8 \block[9].zbuf_pg_ena_I.genblk1.cell0_I  (.A(\block[9].l_ena ),
    .X(\block[9].zbuf_pg_ena_I.z ));
 sg13g2_buf_2 \branch_addr_match_buf_I[0].genblk1.cell0_I  (.A(spine_iw[7]),
    .X(\branch_addr_match_buf_I[0].z ));
 sg13g2_buf_2 \branch_addr_match_buf_I[1].genblk1.cell0_I  (.A(spine_iw[8]),
    .X(\branch_addr_match_buf_I[1].z ));
 sg13g2_buf_2 \branch_addr_match_buf_I[2].genblk1.cell0_I  (.A(spine_iw[9]),
    .X(\branch_addr_match_buf_I[2].z ));
 sg13g2_buf_2 \branch_addr_match_buf_I[3].genblk1.cell0_I  (.A(spine_iw[10]),
    .X(\branch_addr_match_buf_I[3].z ));
 sg13g2_buf_2 \branch_ena_buf_I.genblk1.cell0_I  (.A(spine_iw[1]),
    .X(\branch_ena_buf_I.z ));
 sg13g2_buf_8 \branch_sel_buf_I.genblk1.cell0_I  (.A(\branch_sel_buf_I.a ),
    .X(branch_sel));
 sg13g2_inv_2 \branch_sel_n_buf_I.genblk1.cell0_I  (.Y(branch_sel_n),
    .A(branch_sel));
 sg13g2_buf_8 \buf_bus_ena_I.genblk1.cell0_I  (.A(branch_sel),
    .X(\buf_bus_ena_I.z ));
 sg13g2_buf_8 \buf_bus_sel_I[0].genblk1.cell0_I  (.A(spine_iw[2]),
    .X(\block[0].genblk1.mux4_sel_buf_I[0].a ));
 sg13g2_buf_8 \buf_bus_sel_I[1].genblk1.cell0_I  (.A(spine_iw[3]),
    .X(\block[0].genblk1.mux4_sel_buf_I[1].a ));
 sg13g2_buf_8 \buf_bus_sel_I[2].genblk1.cell0_I  (.A(spine_iw[4]),
    .X(\buf_bus_sel_I[2].z ));
 sg13g2_buf_8 \buf_bus_sel_I[3].genblk1.cell0_I  (.A(spine_iw[5]),
    .X(\buf_bus_sel_I[3].z ));
 sg13g2_buf_8 \buf_bus_sel_I[4].genblk1.cell0_I  (.A(spine_iw[6]),
    .X(\buf_bus_sel_I[4].z ));
 sg13g2_buf_2 \buf_spine_ow_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[0].z ),
    .X(\buf_spine_ow_I[0].z ));
 sg13g2_buf_2 \buf_spine_ow_I[10].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[10].z ),
    .X(\buf_spine_ow_I[10].z ));
 sg13g2_buf_2 \buf_spine_ow_I[11].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[11].z ),
    .X(\buf_spine_ow_I[11].z ));
 sg13g2_buf_2 \buf_spine_ow_I[12].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[12].z ),
    .X(\buf_spine_ow_I[12].z ));
 sg13g2_buf_2 \buf_spine_ow_I[13].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[13].z ),
    .X(\buf_spine_ow_I[13].z ));
 sg13g2_buf_2 \buf_spine_ow_I[14].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[14].z ),
    .X(\buf_spine_ow_I[14].z ));
 sg13g2_buf_2 \buf_spine_ow_I[15].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[15].z ),
    .X(\buf_spine_ow_I[15].z ));
 sg13g2_buf_2 \buf_spine_ow_I[16].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[16].z ),
    .X(\buf_spine_ow_I[16].z ));
 sg13g2_buf_2 \buf_spine_ow_I[17].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[17].z ),
    .X(\buf_spine_ow_I[17].z ));
 sg13g2_buf_2 \buf_spine_ow_I[18].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[18].z ),
    .X(\buf_spine_ow_I[18].z ));
 sg13g2_buf_2 \buf_spine_ow_I[19].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[19].z ),
    .X(\buf_spine_ow_I[19].z ));
 sg13g2_buf_2 \buf_spine_ow_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[1].z ),
    .X(\buf_spine_ow_I[1].z ));
 sg13g2_buf_2 \buf_spine_ow_I[20].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[20].z ),
    .X(\buf_spine_ow_I[20].z ));
 sg13g2_buf_2 \buf_spine_ow_I[21].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[21].z ),
    .X(\buf_spine_ow_I[21].z ));
 sg13g2_buf_2 \buf_spine_ow_I[22].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[22].z ),
    .X(\buf_spine_ow_I[22].z ));
 sg13g2_buf_2 \buf_spine_ow_I[23].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[23].z ),
    .X(\buf_spine_ow_I[23].z ));
 sg13g2_buf_2 \buf_spine_ow_I[2].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[2].z ),
    .X(\buf_spine_ow_I[2].z ));
 sg13g2_buf_2 \buf_spine_ow_I[3].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[3].z ),
    .X(\buf_spine_ow_I[3].z ));
 sg13g2_buf_2 \buf_spine_ow_I[4].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[4].z ),
    .X(\buf_spine_ow_I[4].z ));
 sg13g2_buf_2 \buf_spine_ow_I[5].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[5].z ),
    .X(\buf_spine_ow_I[5].z ));
 sg13g2_buf_2 \buf_spine_ow_I[6].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[6].z ),
    .X(\buf_spine_ow_I[6].z ));
 sg13g2_buf_2 \buf_spine_ow_I[7].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[7].z ),
    .X(\buf_spine_ow_I[7].z ));
 sg13g2_buf_2 \buf_spine_ow_I[8].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[8].z ),
    .X(\buf_spine_ow_I[8].z ));
 sg13g2_buf_2 \buf_spine_ow_I[9].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[9].z ),
    .X(\buf_spine_ow_I[9].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[0].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[10].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[11].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[12].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[13].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[14].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[15].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[16].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[17].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[18].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[19].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[1].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[20].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[21].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[22].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[23].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[2].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[3].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[4].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[5].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[6].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[7].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[8].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ));
 sg13g2_ebufn_4 \bus_pull_ow_I[9].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(branch_sel_n_tbe),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ));
 sg13g2_tielo \bus_pull_tie_I.genblk1.cell0_I  (.L_LO(\bus_pull_ow_I[0].a ));
 sg13g2_antennanp \diode_spine_I[0].cell0_I  (.A(spine_iw[0]));
 sg13g2_antennanp \diode_spine_I[10].cell0_I  (.A(spine_iw[10]));
 sg13g2_antennanp \diode_spine_I[11].cell0_I  (.A(spine_iw[11]));
 sg13g2_antennanp \diode_spine_I[12].cell0_I  (.A(spine_iw[12]));
 sg13g2_antennanp \diode_spine_I[13].cell0_I  (.A(spine_iw[13]));
 sg13g2_antennanp \diode_spine_I[14].cell0_I  (.A(spine_iw[14]));
 sg13g2_antennanp \diode_spine_I[15].cell0_I  (.A(spine_iw[15]));
 sg13g2_antennanp \diode_spine_I[16].cell0_I  (.A(spine_iw[16]));
 sg13g2_antennanp \diode_spine_I[17].cell0_I  (.A(spine_iw[17]));
 sg13g2_antennanp \diode_spine_I[18].cell0_I  (.A(spine_iw[18]));
 sg13g2_antennanp \diode_spine_I[19].cell0_I  (.A(spine_iw[19]));
 sg13g2_antennanp \diode_spine_I[1].cell0_I  (.A(spine_iw[1]));
 sg13g2_antennanp \diode_spine_I[20].cell0_I  (.A(spine_iw[20]));
 sg13g2_antennanp \diode_spine_I[21].cell0_I  (.A(spine_iw[21]));
 sg13g2_antennanp \diode_spine_I[22].cell0_I  (.A(spine_iw[22]));
 sg13g2_antennanp \diode_spine_I[23].cell0_I  (.A(spine_iw[23]));
 sg13g2_antennanp \diode_spine_I[24].cell0_I  (.A(spine_iw[24]));
 sg13g2_antennanp \diode_spine_I[25].cell0_I  (.A(spine_iw[25]));
 sg13g2_antennanp \diode_spine_I[26].cell0_I  (.A(spine_iw[26]));
 sg13g2_antennanp \diode_spine_I[27].cell0_I  (.A(spine_iw[27]));
 sg13g2_antennanp \diode_spine_I[28].cell0_I  (.A(spine_iw[28]));
 sg13g2_antennanp \diode_spine_I[29].cell0_I  (.A(spine_iw[29]));
 sg13g2_antennanp \diode_spine_I[2].cell0_I  (.A(spine_iw[2]));
 sg13g2_antennanp \diode_spine_I[3].cell0_I  (.A(spine_iw[3]));
 sg13g2_antennanp \diode_spine_I[4].cell0_I  (.A(spine_iw[4]));
 sg13g2_antennanp \diode_spine_I[5].cell0_I  (.A(spine_iw[5]));
 sg13g2_antennanp \diode_spine_I[6].cell0_I  (.A(spine_iw[6]));
 sg13g2_antennanp \diode_spine_I[7].cell0_I  (.A(spine_iw[7]));
 sg13g2_antennanp \diode_spine_I[8].cell0_I  (.A(spine_iw[8]));
 sg13g2_antennanp \diode_spine_I[9].cell0_I  (.A(spine_iw[9]));
 sg13g2_inv_8 \tbuf_row_ena_I.cell0_I  (.Y(branch_sel_tbe),
    .A(branch_sel));
 sg13g2_inv_8 \tbuf_row_ena_n_I.cell0_I  (.Y(branch_sel_n_tbe),
    .A(branch_sel_n));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[0].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[0].z ),
    .A(\buf_spine_ow_I[0].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[10].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[10].z ),
    .A(\buf_spine_ow_I[10].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[11].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[11].z ),
    .A(\buf_spine_ow_I[11].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[12].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[12].z ),
    .A(\buf_spine_ow_I[12].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[13].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[13].z ),
    .A(\buf_spine_ow_I[13].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[14].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[14].z ),
    .A(\buf_spine_ow_I[14].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[15].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[15].z ),
    .A(\buf_spine_ow_I[15].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[16].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[16].z ),
    .A(\buf_spine_ow_I[16].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[17].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[17].z ),
    .A(\buf_spine_ow_I[17].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[18].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[18].z ),
    .A(\buf_spine_ow_I[18].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[19].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[19].z ),
    .A(\buf_spine_ow_I[19].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[1].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[1].z ),
    .A(\buf_spine_ow_I[1].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[20].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[20].z ),
    .A(\buf_spine_ow_I[20].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[21].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[21].z ),
    .A(\buf_spine_ow_I[21].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[22].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[22].z ),
    .A(\buf_spine_ow_I[22].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[23].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[23].z ),
    .A(\buf_spine_ow_I[23].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[2].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[2].z ),
    .A(\buf_spine_ow_I[2].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[3].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[3].z ),
    .A(\buf_spine_ow_I[3].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[4].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[4].z ),
    .A(\buf_spine_ow_I[4].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[5].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[5].z ),
    .A(\buf_spine_ow_I[5].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[6].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[6].z ),
    .A(\buf_spine_ow_I[6].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[7].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[7].z ),
    .A(\buf_spine_ow_I[7].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[8].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[8].z ),
    .A(\buf_spine_ow_I[8].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_ebufn_8 \tbuf_spine_ow_I[9].genblk1.cell0_I  (.Z(\tbuf_spine_ow_I[9].z ),
    .A(\buf_spine_ow_I[9].z ),
    .TE_B(branch_sel_tbe));
 sg13g2_tielo \tie_I.genblk1.cell0_I  (.L_LO(k_zero));
 sg13g2_tiehi \tie_I.genblk2.cell1_I  (.L_HI(k_one));
 sg13g2_tielo \tie_spine_guard_I[0].genblk1.cell0_I  (.L_LO(so_gl));
 sg13g2_tielo \tie_spine_guard_I[1].genblk1.cell0_I  (.L_LO(so_gh));
 sg13g2_and2_2 \zbuf_bus_iw_I[0].genblk1.cell0_I  (.A(spine_iw[11]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[0].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[0].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[0].genblk1.l ),
    .X(\block[0].zbuf_iw_I[0].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[10].genblk1.cell0_I  (.A(spine_iw[21]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[10].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[10].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[10].genblk1.l ),
    .X(\block[0].zbuf_iw_I[10].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[11].genblk1.cell0_I  (.A(spine_iw[22]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[11].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[11].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[11].genblk1.l ),
    .X(\block[0].zbuf_iw_I[11].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[12].genblk1.cell0_I  (.A(spine_iw[23]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[12].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[12].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[12].genblk1.l ),
    .X(\block[0].zbuf_iw_I[12].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[13].genblk1.cell0_I  (.A(spine_iw[24]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[13].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[13].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[13].genblk1.l ),
    .X(\block[0].zbuf_iw_I[13].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[14].genblk1.cell0_I  (.A(spine_iw[25]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[14].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[14].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[14].genblk1.l ),
    .X(\block[0].zbuf_iw_I[14].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[15].genblk1.cell0_I  (.A(spine_iw[26]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[15].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[15].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[15].genblk1.l ),
    .X(\block[0].zbuf_iw_I[15].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[16].genblk1.cell0_I  (.A(spine_iw[27]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[16].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[16].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[16].genblk1.l ),
    .X(\block[0].zbuf_iw_I[16].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[17].genblk1.cell0_I  (.A(spine_iw[28]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[17].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[17].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[17].genblk1.l ),
    .X(\block[0].zbuf_iw_I[17].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[1].genblk1.cell0_I  (.A(spine_iw[12]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[1].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[1].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[1].genblk1.l ),
    .X(\block[0].zbuf_iw_I[1].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[2].genblk1.cell0_I  (.A(spine_iw[13]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[2].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[2].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[2].genblk1.l ),
    .X(\block[0].zbuf_iw_I[2].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[3].genblk1.cell0_I  (.A(spine_iw[14]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[3].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[3].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[3].genblk1.l ),
    .X(\block[0].zbuf_iw_I[3].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[4].genblk1.cell0_I  (.A(spine_iw[15]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[4].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[4].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[4].genblk1.l ),
    .X(\block[0].zbuf_iw_I[4].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[5].genblk1.cell0_I  (.A(spine_iw[16]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[5].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[5].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[5].genblk1.l ),
    .X(\block[0].zbuf_iw_I[5].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[6].genblk1.cell0_I  (.A(spine_iw[17]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[6].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[6].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[6].genblk1.l ),
    .X(\block[0].zbuf_iw_I[6].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[7].genblk1.cell0_I  (.A(spine_iw[18]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[7].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[7].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[7].genblk1.l ),
    .X(\block[0].zbuf_iw_I[7].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[8].genblk1.cell0_I  (.A(spine_iw[19]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[8].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[8].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[8].genblk1.l ),
    .X(\block[0].zbuf_iw_I[8].a ));
 sg13g2_and2_2 \zbuf_bus_iw_I[9].genblk1.cell0_I  (.A(spine_iw[20]),
    .B(branch_sel),
    .X(\zbuf_bus_iw_I[9].genblk1.l ));
 sg13g2_buf_8 \zbuf_bus_iw_I[9].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[9].genblk1.l ),
    .X(\block[0].zbuf_iw_I[9].a ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_fill_2 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_414 ();
 sg13g2_decap_8 FILLER_0_421 ();
 sg13g2_decap_8 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_0_435 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_decap_8 FILLER_0_449 ();
 sg13g2_decap_8 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_463 ();
 sg13g2_decap_8 FILLER_0_470 ();
 sg13g2_decap_8 FILLER_0_477 ();
 sg13g2_decap_8 FILLER_0_484 ();
 sg13g2_decap_8 FILLER_0_491 ();
 sg13g2_decap_8 FILLER_0_498 ();
 sg13g2_decap_8 FILLER_0_505 ();
 sg13g2_decap_8 FILLER_0_512 ();
 sg13g2_decap_4 FILLER_0_519 ();
 sg13g2_fill_2 FILLER_0_523 ();
 sg13g2_decap_8 FILLER_0_528 ();
 sg13g2_decap_8 FILLER_0_535 ();
 sg13g2_decap_8 FILLER_0_542 ();
 sg13g2_decap_8 FILLER_0_549 ();
 sg13g2_decap_8 FILLER_0_556 ();
 sg13g2_decap_8 FILLER_0_563 ();
 sg13g2_decap_8 FILLER_0_570 ();
 sg13g2_decap_8 FILLER_0_577 ();
 sg13g2_decap_8 FILLER_0_584 ();
 sg13g2_decap_8 FILLER_0_591 ();
 sg13g2_decap_8 FILLER_0_598 ();
 sg13g2_decap_8 FILLER_0_605 ();
 sg13g2_decap_8 FILLER_0_612 ();
 sg13g2_decap_8 FILLER_0_619 ();
 sg13g2_decap_8 FILLER_0_626 ();
 sg13g2_decap_8 FILLER_0_633 ();
 sg13g2_decap_8 FILLER_0_640 ();
 sg13g2_decap_8 FILLER_0_647 ();
 sg13g2_decap_8 FILLER_0_654 ();
 sg13g2_decap_8 FILLER_0_661 ();
 sg13g2_decap_8 FILLER_0_668 ();
 sg13g2_decap_8 FILLER_0_675 ();
 sg13g2_decap_8 FILLER_0_682 ();
 sg13g2_decap_8 FILLER_0_689 ();
 sg13g2_decap_8 FILLER_0_696 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_787 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_899 ();
 sg13g2_decap_8 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_913 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_8 FILLER_0_1025 ();
 sg13g2_decap_8 FILLER_0_1032 ();
 sg13g2_decap_8 FILLER_0_1039 ();
 sg13g2_decap_8 FILLER_0_1046 ();
 sg13g2_decap_8 FILLER_0_1053 ();
 sg13g2_decap_8 FILLER_0_1060 ();
 sg13g2_decap_8 FILLER_0_1067 ();
 sg13g2_decap_8 FILLER_0_1074 ();
 sg13g2_decap_8 FILLER_0_1081 ();
 sg13g2_decap_8 FILLER_0_1088 ();
 sg13g2_decap_8 FILLER_0_1095 ();
 sg13g2_decap_8 FILLER_0_1102 ();
 sg13g2_decap_8 FILLER_0_1109 ();
 sg13g2_decap_8 FILLER_0_1116 ();
 sg13g2_decap_8 FILLER_0_1123 ();
 sg13g2_decap_8 FILLER_0_1130 ();
 sg13g2_decap_8 FILLER_0_1137 ();
 sg13g2_decap_8 FILLER_0_1144 ();
 sg13g2_decap_8 FILLER_0_1151 ();
 sg13g2_decap_8 FILLER_0_1158 ();
 sg13g2_decap_8 FILLER_0_1165 ();
 sg13g2_decap_8 FILLER_0_1172 ();
 sg13g2_decap_8 FILLER_0_1179 ();
 sg13g2_decap_8 FILLER_0_1186 ();
 sg13g2_decap_8 FILLER_0_1193 ();
 sg13g2_decap_8 FILLER_0_1200 ();
 sg13g2_decap_8 FILLER_0_1207 ();
 sg13g2_decap_8 FILLER_0_1214 ();
 sg13g2_decap_8 FILLER_0_1221 ();
 sg13g2_decap_8 FILLER_0_1228 ();
 sg13g2_fill_2 FILLER_0_1235 ();
 sg13g2_fill_1 FILLER_0_1237 ();
 sg13g2_decap_8 FILLER_0_1241 ();
 sg13g2_decap_8 FILLER_0_1248 ();
 sg13g2_decap_8 FILLER_0_1255 ();
 sg13g2_decap_8 FILLER_0_1262 ();
 sg13g2_decap_8 FILLER_0_1269 ();
 sg13g2_decap_8 FILLER_0_1276 ();
 sg13g2_decap_8 FILLER_0_1283 ();
 sg13g2_decap_8 FILLER_0_1290 ();
 sg13g2_decap_8 FILLER_0_1297 ();
 sg13g2_decap_8 FILLER_0_1304 ();
 sg13g2_decap_8 FILLER_0_1311 ();
 sg13g2_decap_8 FILLER_0_1318 ();
 sg13g2_decap_8 FILLER_0_1325 ();
 sg13g2_decap_8 FILLER_0_1332 ();
 sg13g2_decap_8 FILLER_0_1339 ();
 sg13g2_decap_8 FILLER_0_1346 ();
 sg13g2_decap_8 FILLER_0_1353 ();
 sg13g2_decap_8 FILLER_0_1360 ();
 sg13g2_decap_8 FILLER_0_1367 ();
 sg13g2_decap_8 FILLER_0_1374 ();
 sg13g2_decap_8 FILLER_0_1381 ();
 sg13g2_decap_8 FILLER_0_1388 ();
 sg13g2_decap_8 FILLER_0_1395 ();
 sg13g2_decap_8 FILLER_0_1402 ();
 sg13g2_decap_8 FILLER_0_1409 ();
 sg13g2_decap_8 FILLER_0_1416 ();
 sg13g2_decap_8 FILLER_0_1423 ();
 sg13g2_decap_8 FILLER_0_1430 ();
 sg13g2_decap_8 FILLER_0_1437 ();
 sg13g2_decap_8 FILLER_0_1444 ();
 sg13g2_decap_8 FILLER_0_1451 ();
 sg13g2_decap_8 FILLER_0_1458 ();
 sg13g2_decap_8 FILLER_0_1465 ();
 sg13g2_decap_8 FILLER_0_1472 ();
 sg13g2_decap_8 FILLER_0_1479 ();
 sg13g2_decap_8 FILLER_0_1486 ();
 sg13g2_decap_8 FILLER_0_1493 ();
 sg13g2_decap_8 FILLER_0_1500 ();
 sg13g2_decap_8 FILLER_0_1507 ();
 sg13g2_decap_8 FILLER_0_1514 ();
 sg13g2_decap_8 FILLER_0_1521 ();
 sg13g2_decap_8 FILLER_0_1528 ();
 sg13g2_decap_8 FILLER_0_1535 ();
 sg13g2_decap_8 FILLER_0_1542 ();
 sg13g2_decap_8 FILLER_0_1549 ();
 sg13g2_decap_8 FILLER_0_1556 ();
 sg13g2_decap_8 FILLER_0_1563 ();
 sg13g2_decap_8 FILLER_0_1570 ();
 sg13g2_decap_8 FILLER_0_1577 ();
 sg13g2_decap_8 FILLER_0_1584 ();
 sg13g2_decap_8 FILLER_0_1591 ();
 sg13g2_decap_8 FILLER_0_1598 ();
 sg13g2_decap_8 FILLER_0_1605 ();
 sg13g2_decap_8 FILLER_0_1612 ();
 sg13g2_decap_8 FILLER_0_1619 ();
 sg13g2_decap_8 FILLER_0_1626 ();
 sg13g2_decap_8 FILLER_0_1633 ();
 sg13g2_decap_8 FILLER_0_1640 ();
 sg13g2_decap_8 FILLER_0_1647 ();
 sg13g2_decap_8 FILLER_0_1654 ();
 sg13g2_decap_8 FILLER_0_1661 ();
 sg13g2_decap_8 FILLER_0_1668 ();
 sg13g2_decap_8 FILLER_0_1675 ();
 sg13g2_decap_8 FILLER_0_1682 ();
 sg13g2_decap_8 FILLER_0_1689 ();
 sg13g2_decap_8 FILLER_0_1696 ();
 sg13g2_decap_8 FILLER_0_1703 ();
 sg13g2_decap_8 FILLER_0_1710 ();
 sg13g2_decap_8 FILLER_0_1717 ();
 sg13g2_decap_8 FILLER_0_1724 ();
 sg13g2_decap_8 FILLER_0_1731 ();
 sg13g2_decap_8 FILLER_0_1738 ();
 sg13g2_decap_8 FILLER_0_1745 ();
 sg13g2_decap_8 FILLER_0_1752 ();
 sg13g2_decap_8 FILLER_0_1759 ();
 sg13g2_decap_8 FILLER_0_1766 ();
 sg13g2_decap_8 FILLER_0_1773 ();
 sg13g2_decap_8 FILLER_0_1780 ();
 sg13g2_decap_8 FILLER_0_1787 ();
 sg13g2_decap_8 FILLER_0_1794 ();
 sg13g2_decap_8 FILLER_0_1801 ();
 sg13g2_decap_8 FILLER_0_1808 ();
 sg13g2_decap_8 FILLER_0_1815 ();
 sg13g2_decap_8 FILLER_0_1822 ();
 sg13g2_decap_8 FILLER_0_1829 ();
 sg13g2_decap_8 FILLER_0_1836 ();
 sg13g2_decap_8 FILLER_0_1843 ();
 sg13g2_decap_8 FILLER_0_1850 ();
 sg13g2_decap_8 FILLER_0_1857 ();
 sg13g2_decap_8 FILLER_0_1864 ();
 sg13g2_decap_8 FILLER_0_1871 ();
 sg13g2_decap_8 FILLER_0_1878 ();
 sg13g2_decap_8 FILLER_0_1885 ();
 sg13g2_decap_8 FILLER_0_1892 ();
 sg13g2_decap_8 FILLER_0_1899 ();
 sg13g2_decap_8 FILLER_0_1906 ();
 sg13g2_fill_2 FILLER_0_1913 ();
 sg13g2_fill_1 FILLER_0_1915 ();
 sg13g2_decap_8 FILLER_0_1919 ();
 sg13g2_decap_8 FILLER_0_1926 ();
 sg13g2_decap_8 FILLER_0_1933 ();
 sg13g2_decap_8 FILLER_0_1940 ();
 sg13g2_decap_8 FILLER_0_1947 ();
 sg13g2_decap_8 FILLER_0_1954 ();
 sg13g2_decap_8 FILLER_0_1961 ();
 sg13g2_decap_8 FILLER_0_1968 ();
 sg13g2_decap_8 FILLER_0_1975 ();
 sg13g2_decap_8 FILLER_0_1982 ();
 sg13g2_decap_8 FILLER_0_1989 ();
 sg13g2_decap_8 FILLER_0_1996 ();
 sg13g2_decap_8 FILLER_0_2003 ();
 sg13g2_decap_8 FILLER_0_2010 ();
 sg13g2_decap_8 FILLER_0_2017 ();
 sg13g2_decap_8 FILLER_0_2024 ();
 sg13g2_decap_8 FILLER_0_2031 ();
 sg13g2_decap_8 FILLER_0_2038 ();
 sg13g2_decap_8 FILLER_0_2045 ();
 sg13g2_decap_8 FILLER_0_2052 ();
 sg13g2_decap_8 FILLER_0_2059 ();
 sg13g2_decap_8 FILLER_0_2066 ();
 sg13g2_decap_8 FILLER_0_2073 ();
 sg13g2_decap_8 FILLER_0_2080 ();
 sg13g2_decap_8 FILLER_0_2087 ();
 sg13g2_decap_4 FILLER_0_2094 ();
 sg13g2_fill_2 FILLER_0_2098 ();
 sg13g2_decap_8 FILLER_0_2103 ();
 sg13g2_decap_8 FILLER_0_2110 ();
 sg13g2_decap_8 FILLER_0_2117 ();
 sg13g2_decap_8 FILLER_0_2124 ();
 sg13g2_decap_8 FILLER_0_2131 ();
 sg13g2_decap_8 FILLER_0_2138 ();
 sg13g2_decap_8 FILLER_0_2145 ();
 sg13g2_decap_8 FILLER_0_2155 ();
 sg13g2_decap_8 FILLER_0_2162 ();
 sg13g2_fill_2 FILLER_0_2169 ();
 sg13g2_fill_1 FILLER_0_2171 ();
 sg13g2_decap_8 FILLER_0_2175 ();
 sg13g2_decap_8 FILLER_0_2182 ();
 sg13g2_decap_8 FILLER_0_2189 ();
 sg13g2_decap_8 FILLER_0_2196 ();
 sg13g2_decap_8 FILLER_0_2203 ();
 sg13g2_decap_4 FILLER_0_2210 ();
 sg13g2_fill_1 FILLER_0_2214 ();
 sg13g2_decap_8 FILLER_0_2218 ();
 sg13g2_decap_8 FILLER_0_2225 ();
 sg13g2_decap_8 FILLER_0_2232 ();
 sg13g2_decap_8 FILLER_0_2239 ();
 sg13g2_decap_8 FILLER_0_2246 ();
 sg13g2_decap_8 FILLER_0_2253 ();
 sg13g2_decap_8 FILLER_0_2260 ();
 sg13g2_decap_8 FILLER_0_2267 ();
 sg13g2_decap_8 FILLER_0_2274 ();
 sg13g2_decap_8 FILLER_0_2281 ();
 sg13g2_decap_8 FILLER_0_2288 ();
 sg13g2_decap_8 FILLER_0_2295 ();
 sg13g2_decap_8 FILLER_0_2302 ();
 sg13g2_decap_8 FILLER_0_2309 ();
 sg13g2_decap_8 FILLER_0_2316 ();
 sg13g2_decap_8 FILLER_0_2323 ();
 sg13g2_decap_8 FILLER_0_2330 ();
 sg13g2_decap_8 FILLER_0_2337 ();
 sg13g2_decap_8 FILLER_0_2344 ();
 sg13g2_decap_8 FILLER_0_2351 ();
 sg13g2_decap_8 FILLER_0_2358 ();
 sg13g2_decap_8 FILLER_0_2365 ();
 sg13g2_decap_8 FILLER_0_2372 ();
 sg13g2_decap_8 FILLER_0_2379 ();
 sg13g2_decap_8 FILLER_0_2386 ();
 sg13g2_decap_8 FILLER_0_2393 ();
 sg13g2_decap_8 FILLER_0_2400 ();
 sg13g2_decap_8 FILLER_0_2407 ();
 sg13g2_decap_8 FILLER_0_2414 ();
 sg13g2_decap_8 FILLER_0_2421 ();
 sg13g2_decap_8 FILLER_0_2428 ();
 sg13g2_decap_8 FILLER_0_2435 ();
 sg13g2_decap_8 FILLER_0_2442 ();
 sg13g2_decap_8 FILLER_0_2449 ();
 sg13g2_decap_8 FILLER_0_2456 ();
 sg13g2_decap_8 FILLER_0_2463 ();
 sg13g2_decap_8 FILLER_0_2470 ();
 sg13g2_decap_8 FILLER_0_2477 ();
 sg13g2_decap_8 FILLER_0_2484 ();
 sg13g2_decap_8 FILLER_0_2491 ();
 sg13g2_decap_8 FILLER_0_2498 ();
 sg13g2_decap_8 FILLER_0_2505 ();
 sg13g2_decap_8 FILLER_0_2512 ();
 sg13g2_decap_8 FILLER_0_2519 ();
 sg13g2_decap_8 FILLER_0_2526 ();
 sg13g2_decap_8 FILLER_0_2533 ();
 sg13g2_decap_8 FILLER_0_2540 ();
 sg13g2_decap_8 FILLER_0_2547 ();
 sg13g2_decap_8 FILLER_0_2554 ();
 sg13g2_decap_8 FILLER_0_2561 ();
 sg13g2_decap_8 FILLER_0_2568 ();
 sg13g2_decap_8 FILLER_0_2575 ();
 sg13g2_decap_8 FILLER_0_2582 ();
 sg13g2_decap_8 FILLER_0_2589 ();
 sg13g2_decap_8 FILLER_0_2596 ();
 sg13g2_decap_8 FILLER_0_2603 ();
 sg13g2_decap_8 FILLER_0_2610 ();
 sg13g2_decap_8 FILLER_0_2617 ();
 sg13g2_decap_8 FILLER_0_2624 ();
 sg13g2_decap_8 FILLER_0_2631 ();
 sg13g2_decap_8 FILLER_0_2638 ();
 sg13g2_decap_8 FILLER_0_2645 ();
 sg13g2_decap_8 FILLER_0_2652 ();
 sg13g2_decap_8 FILLER_0_2659 ();
 sg13g2_decap_8 FILLER_0_2666 ();
 sg13g2_decap_8 FILLER_0_2673 ();
 sg13g2_decap_8 FILLER_0_2680 ();
 sg13g2_decap_8 FILLER_0_2687 ();
 sg13g2_decap_4 FILLER_0_2694 ();
 sg13g2_fill_2 FILLER_0_2698 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_fill_1 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_75 ();
 sg13g2_decap_8 FILLER_1_82 ();
 sg13g2_decap_8 FILLER_1_89 ();
 sg13g2_decap_8 FILLER_1_96 ();
 sg13g2_decap_8 FILLER_1_103 ();
 sg13g2_decap_8 FILLER_1_110 ();
 sg13g2_decap_8 FILLER_1_117 ();
 sg13g2_decap_8 FILLER_1_124 ();
 sg13g2_decap_8 FILLER_1_131 ();
 sg13g2_decap_8 FILLER_1_138 ();
 sg13g2_decap_8 FILLER_1_145 ();
 sg13g2_decap_8 FILLER_1_152 ();
 sg13g2_decap_8 FILLER_1_159 ();
 sg13g2_decap_8 FILLER_1_166 ();
 sg13g2_decap_8 FILLER_1_173 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_208 ();
 sg13g2_decap_8 FILLER_1_215 ();
 sg13g2_decap_8 FILLER_1_222 ();
 sg13g2_decap_8 FILLER_1_229 ();
 sg13g2_decap_8 FILLER_1_236 ();
 sg13g2_decap_8 FILLER_1_243 ();
 sg13g2_decap_8 FILLER_1_250 ();
 sg13g2_decap_8 FILLER_1_257 ();
 sg13g2_fill_2 FILLER_1_264 ();
 sg13g2_fill_1 FILLER_1_266 ();
 sg13g2_fill_2 FILLER_1_280 ();
 sg13g2_fill_2 FILLER_1_288 ();
 sg13g2_fill_2 FILLER_1_296 ();
 sg13g2_fill_2 FILLER_1_304 ();
 sg13g2_fill_2 FILLER_1_312 ();
 sg13g2_fill_2 FILLER_1_320 ();
 sg13g2_fill_2 FILLER_1_328 ();
 sg13g2_fill_2 FILLER_1_336 ();
 sg13g2_fill_2 FILLER_1_344 ();
 sg13g2_fill_2 FILLER_1_352 ();
 sg13g2_fill_2 FILLER_1_360 ();
 sg13g2_fill_2 FILLER_1_368 ();
 sg13g2_fill_2 FILLER_1_376 ();
 sg13g2_fill_2 FILLER_1_384 ();
 sg13g2_fill_2 FILLER_1_392 ();
 sg13g2_fill_2 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_decap_8 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_1_435 ();
 sg13g2_decap_8 FILLER_1_442 ();
 sg13g2_decap_8 FILLER_1_449 ();
 sg13g2_decap_8 FILLER_1_456 ();
 sg13g2_decap_8 FILLER_1_463 ();
 sg13g2_decap_8 FILLER_1_470 ();
 sg13g2_decap_8 FILLER_1_477 ();
 sg13g2_decap_8 FILLER_1_484 ();
 sg13g2_decap_8 FILLER_1_491 ();
 sg13g2_decap_8 FILLER_1_498 ();
 sg13g2_decap_8 FILLER_1_505 ();
 sg13g2_decap_8 FILLER_1_512 ();
 sg13g2_fill_1 FILLER_1_519 ();
 sg13g2_fill_2 FILLER_1_527 ();
 sg13g2_fill_1 FILLER_1_535 ();
 sg13g2_decap_4 FILLER_1_539 ();
 sg13g2_fill_1 FILLER_1_543 ();
 sg13g2_decap_4 FILLER_1_547 ();
 sg13g2_fill_1 FILLER_1_551 ();
 sg13g2_fill_1 FILLER_1_561 ();
 sg13g2_fill_1 FILLER_1_565 ();
 sg13g2_fill_2 FILLER_1_569 ();
 sg13g2_fill_1 FILLER_1_574 ();
 sg13g2_fill_1 FILLER_1_578 ();
 sg13g2_fill_2 FILLER_1_585 ();
 sg13g2_fill_1 FILLER_1_587 ();
 sg13g2_decap_4 FILLER_1_591 ();
 sg13g2_fill_2 FILLER_1_607 ();
 sg13g2_fill_1 FILLER_1_618 ();
 sg13g2_fill_2 FILLER_1_625 ();
 sg13g2_decap_4 FILLER_1_639 ();
 sg13g2_fill_1 FILLER_1_649 ();
 sg13g2_decap_4 FILLER_1_662 ();
 sg13g2_decap_4 FILLER_1_672 ();
 sg13g2_fill_2 FILLER_1_682 ();
 sg13g2_fill_1 FILLER_1_684 ();
 sg13g2_fill_2 FILLER_1_694 ();
 sg13g2_fill_1 FILLER_1_696 ();
 sg13g2_decap_4 FILLER_1_703 ();
 sg13g2_fill_1 FILLER_1_707 ();
 sg13g2_fill_1 FILLER_1_711 ();
 sg13g2_fill_1 FILLER_1_737 ();
 sg13g2_fill_2 FILLER_1_744 ();
 sg13g2_fill_1 FILLER_1_746 ();
 sg13g2_fill_2 FILLER_1_753 ();
 sg13g2_fill_2 FILLER_1_761 ();
 sg13g2_fill_1 FILLER_1_763 ();
 sg13g2_fill_2 FILLER_1_770 ();
 sg13g2_fill_1 FILLER_1_778 ();
 sg13g2_fill_1 FILLER_1_785 ();
 sg13g2_fill_2 FILLER_1_792 ();
 sg13g2_fill_2 FILLER_1_800 ();
 sg13g2_fill_1 FILLER_1_802 ();
 sg13g2_fill_2 FILLER_1_809 ();
 sg13g2_fill_2 FILLER_1_817 ();
 sg13g2_fill_2 FILLER_1_825 ();
 sg13g2_fill_1 FILLER_1_833 ();
 sg13g2_fill_2 FILLER_1_840 ();
 sg13g2_fill_2 FILLER_1_848 ();
 sg13g2_fill_1 FILLER_1_850 ();
 sg13g2_fill_2 FILLER_1_857 ();
 sg13g2_decap_4 FILLER_1_865 ();
 sg13g2_decap_8 FILLER_1_874 ();
 sg13g2_decap_8 FILLER_1_881 ();
 sg13g2_decap_8 FILLER_1_888 ();
 sg13g2_decap_8 FILLER_1_895 ();
 sg13g2_decap_8 FILLER_1_902 ();
 sg13g2_decap_8 FILLER_1_909 ();
 sg13g2_decap_8 FILLER_1_916 ();
 sg13g2_decap_8 FILLER_1_923 ();
 sg13g2_decap_8 FILLER_1_930 ();
 sg13g2_decap_8 FILLER_1_937 ();
 sg13g2_decap_8 FILLER_1_944 ();
 sg13g2_decap_8 FILLER_1_951 ();
 sg13g2_decap_8 FILLER_1_958 ();
 sg13g2_decap_8 FILLER_1_965 ();
 sg13g2_decap_4 FILLER_1_972 ();
 sg13g2_fill_1 FILLER_1_976 ();
 sg13g2_decap_8 FILLER_1_981 ();
 sg13g2_decap_4 FILLER_1_988 ();
 sg13g2_decap_8 FILLER_1_995 ();
 sg13g2_fill_1 FILLER_1_1005 ();
 sg13g2_fill_1 FILLER_1_1033 ();
 sg13g2_decap_8 FILLER_1_1037 ();
 sg13g2_decap_4 FILLER_1_1044 ();
 sg13g2_decap_8 FILLER_1_1075 ();
 sg13g2_fill_1 FILLER_1_1082 ();
 sg13g2_decap_8 FILLER_1_1086 ();
 sg13g2_fill_2 FILLER_1_1093 ();
 sg13g2_decap_4 FILLER_1_1101 ();
 sg13g2_decap_8 FILLER_1_1108 ();
 sg13g2_fill_2 FILLER_1_1115 ();
 sg13g2_fill_1 FILLER_1_1117 ();
 sg13g2_decap_8 FILLER_1_1121 ();
 sg13g2_fill_2 FILLER_1_1128 ();
 sg13g2_decap_4 FILLER_1_1136 ();
 sg13g2_fill_1 FILLER_1_1140 ();
 sg13g2_decap_4 FILLER_1_1154 ();
 sg13g2_fill_1 FILLER_1_1158 ();
 sg13g2_decap_4 FILLER_1_1162 ();
 sg13g2_fill_2 FILLER_1_1166 ();
 sg13g2_fill_2 FILLER_1_1171 ();
 sg13g2_fill_2 FILLER_1_1182 ();
 sg13g2_fill_2 FILLER_1_1190 ();
 sg13g2_fill_2 FILLER_1_1207 ();
 sg13g2_fill_2 FILLER_1_1215 ();
 sg13g2_fill_1 FILLER_1_1223 ();
 sg13g2_fill_1 FILLER_1_1230 ();
 sg13g2_fill_2 FILLER_1_1237 ();
 sg13g2_fill_2 FILLER_1_1245 ();
 sg13g2_fill_2 FILLER_1_1262 ();
 sg13g2_fill_2 FILLER_1_1270 ();
 sg13g2_fill_2 FILLER_1_1278 ();
 sg13g2_fill_2 FILLER_1_1295 ();
 sg13g2_fill_2 FILLER_1_1321 ();
 sg13g2_fill_1 FILLER_1_1323 ();
 sg13g2_decap_8 FILLER_1_1332 ();
 sg13g2_decap_8 FILLER_1_1339 ();
 sg13g2_decap_8 FILLER_1_1346 ();
 sg13g2_decap_8 FILLER_1_1353 ();
 sg13g2_decap_8 FILLER_1_1360 ();
 sg13g2_decap_8 FILLER_1_1367 ();
 sg13g2_decap_8 FILLER_1_1374 ();
 sg13g2_decap_8 FILLER_1_1381 ();
 sg13g2_decap_8 FILLER_1_1388 ();
 sg13g2_decap_8 FILLER_1_1398 ();
 sg13g2_decap_8 FILLER_1_1405 ();
 sg13g2_decap_8 FILLER_1_1412 ();
 sg13g2_decap_8 FILLER_1_1419 ();
 sg13g2_decap_4 FILLER_1_1426 ();
 sg13g2_fill_2 FILLER_1_1434 ();
 sg13g2_decap_4 FILLER_1_1439 ();
 sg13g2_fill_1 FILLER_1_1443 ();
 sg13g2_decap_4 FILLER_1_1447 ();
 sg13g2_fill_2 FILLER_1_1451 ();
 sg13g2_decap_8 FILLER_1_1456 ();
 sg13g2_decap_8 FILLER_1_1463 ();
 sg13g2_decap_8 FILLER_1_1470 ();
 sg13g2_decap_8 FILLER_1_1480 ();
 sg13g2_decap_4 FILLER_1_1487 ();
 sg13g2_fill_1 FILLER_1_1491 ();
 sg13g2_decap_8 FILLER_1_1495 ();
 sg13g2_decap_8 FILLER_1_1502 ();
 sg13g2_decap_8 FILLER_1_1509 ();
 sg13g2_decap_8 FILLER_1_1516 ();
 sg13g2_decap_8 FILLER_1_1523 ();
 sg13g2_fill_2 FILLER_1_1530 ();
 sg13g2_fill_1 FILLER_1_1532 ();
 sg13g2_decap_4 FILLER_1_1536 ();
 sg13g2_fill_1 FILLER_1_1540 ();
 sg13g2_decap_4 FILLER_1_1544 ();
 sg13g2_fill_1 FILLER_1_1548 ();
 sg13g2_decap_8 FILLER_1_1552 ();
 sg13g2_decap_8 FILLER_1_1559 ();
 sg13g2_decap_4 FILLER_1_1569 ();
 sg13g2_fill_1 FILLER_1_1573 ();
 sg13g2_decap_4 FILLER_1_1577 ();
 sg13g2_decap_4 FILLER_1_1584 ();
 sg13g2_fill_1 FILLER_1_1588 ();
 sg13g2_decap_8 FILLER_1_1592 ();
 sg13g2_decap_8 FILLER_1_1599 ();
 sg13g2_decap_8 FILLER_1_1606 ();
 sg13g2_decap_8 FILLER_1_1613 ();
 sg13g2_fill_1 FILLER_1_1620 ();
 sg13g2_fill_2 FILLER_1_1652 ();
 sg13g2_fill_2 FILLER_1_1660 ();
 sg13g2_fill_1 FILLER_1_1668 ();
 sg13g2_fill_2 FILLER_1_1675 ();
 sg13g2_fill_2 FILLER_1_1683 ();
 sg13g2_fill_2 FILLER_1_1691 ();
 sg13g2_fill_2 FILLER_1_1699 ();
 sg13g2_fill_2 FILLER_1_1707 ();
 sg13g2_fill_2 FILLER_1_1715 ();
 sg13g2_fill_2 FILLER_1_1723 ();
 sg13g2_fill_1 FILLER_1_1725 ();
 sg13g2_fill_2 FILLER_1_1732 ();
 sg13g2_fill_2 FILLER_1_1740 ();
 sg13g2_fill_1 FILLER_1_1748 ();
 sg13g2_fill_2 FILLER_1_1755 ();
 sg13g2_decap_8 FILLER_1_1774 ();
 sg13g2_decap_8 FILLER_1_1781 ();
 sg13g2_decap_8 FILLER_1_1788 ();
 sg13g2_decap_8 FILLER_1_1795 ();
 sg13g2_decap_4 FILLER_1_1802 ();
 sg13g2_fill_2 FILLER_1_1806 ();
 sg13g2_decap_8 FILLER_1_1821 ();
 sg13g2_decap_8 FILLER_1_1828 ();
 sg13g2_decap_8 FILLER_1_1835 ();
 sg13g2_decap_8 FILLER_1_1842 ();
 sg13g2_decap_8 FILLER_1_1849 ();
 sg13g2_decap_8 FILLER_1_1856 ();
 sg13g2_decap_8 FILLER_1_1863 ();
 sg13g2_decap_8 FILLER_1_1870 ();
 sg13g2_decap_4 FILLER_1_1877 ();
 sg13g2_fill_1 FILLER_1_1881 ();
 sg13g2_decap_8 FILLER_1_1886 ();
 sg13g2_decap_8 FILLER_1_1893 ();
 sg13g2_fill_2 FILLER_1_1903 ();
 sg13g2_fill_1 FILLER_1_1905 ();
 sg13g2_fill_2 FILLER_1_1930 ();
 sg13g2_decap_4 FILLER_1_1935 ();
 sg13g2_fill_1 FILLER_1_1939 ();
 sg13g2_decap_8 FILLER_1_1943 ();
 sg13g2_decap_8 FILLER_1_1950 ();
 sg13g2_fill_2 FILLER_1_1957 ();
 sg13g2_fill_1 FILLER_1_1959 ();
 sg13g2_decap_8 FILLER_1_1963 ();
 sg13g2_fill_2 FILLER_1_1970 ();
 sg13g2_fill_1 FILLER_1_1972 ();
 sg13g2_decap_8 FILLER_1_1976 ();
 sg13g2_fill_2 FILLER_1_1989 ();
 sg13g2_fill_1 FILLER_1_1991 ();
 sg13g2_decap_8 FILLER_1_1995 ();
 sg13g2_decap_8 FILLER_1_2005 ();
 sg13g2_decap_8 FILLER_1_2018 ();
 sg13g2_fill_2 FILLER_1_2025 ();
 sg13g2_fill_2 FILLER_1_2030 ();
 sg13g2_fill_1 FILLER_1_2035 ();
 sg13g2_decap_8 FILLER_1_2042 ();
 sg13g2_decap_8 FILLER_1_2049 ();
 sg13g2_decap_8 FILLER_1_2056 ();
 sg13g2_fill_1 FILLER_1_2063 ();
 sg13g2_fill_1 FILLER_1_2073 ();
 sg13g2_fill_1 FILLER_1_2080 ();
 sg13g2_decap_4 FILLER_1_2087 ();
 sg13g2_fill_2 FILLER_1_2097 ();
 sg13g2_fill_1 FILLER_1_2105 ();
 sg13g2_fill_1 FILLER_1_2112 ();
 sg13g2_fill_2 FILLER_1_2119 ();
 sg13g2_fill_2 FILLER_1_2127 ();
 sg13g2_fill_1 FILLER_1_2144 ();
 sg13g2_fill_2 FILLER_1_2151 ();
 sg13g2_fill_2 FILLER_1_2159 ();
 sg13g2_fill_2 FILLER_1_2167 ();
 sg13g2_fill_2 FILLER_1_2175 ();
 sg13g2_fill_2 FILLER_1_2183 ();
 sg13g2_fill_1 FILLER_1_2185 ();
 sg13g2_fill_1 FILLER_1_2192 ();
 sg13g2_fill_2 FILLER_1_2199 ();
 sg13g2_fill_1 FILLER_1_2201 ();
 sg13g2_fill_1 FILLER_1_2217 ();
 sg13g2_fill_2 FILLER_1_2229 ();
 sg13g2_fill_1 FILLER_1_2231 ();
 sg13g2_decap_8 FILLER_1_2241 ();
 sg13g2_decap_8 FILLER_1_2248 ();
 sg13g2_fill_2 FILLER_1_2255 ();
 sg13g2_fill_1 FILLER_1_2257 ();
 sg13g2_fill_1 FILLER_1_2271 ();
 sg13g2_decap_8 FILLER_1_2287 ();
 sg13g2_decap_8 FILLER_1_2294 ();
 sg13g2_decap_4 FILLER_1_2301 ();
 sg13g2_fill_1 FILLER_1_2305 ();
 sg13g2_decap_8 FILLER_1_2309 ();
 sg13g2_decap_8 FILLER_1_2316 ();
 sg13g2_decap_8 FILLER_1_2323 ();
 sg13g2_fill_2 FILLER_1_2330 ();
 sg13g2_fill_1 FILLER_1_2332 ();
 sg13g2_fill_2 FILLER_1_2340 ();
 sg13g2_decap_4 FILLER_1_2345 ();
 sg13g2_fill_1 FILLER_1_2349 ();
 sg13g2_decap_4 FILLER_1_2353 ();
 sg13g2_fill_2 FILLER_1_2357 ();
 sg13g2_fill_2 FILLER_1_2362 ();
 sg13g2_fill_1 FILLER_1_2364 ();
 sg13g2_decap_4 FILLER_1_2373 ();
 sg13g2_fill_1 FILLER_1_2377 ();
 sg13g2_decap_4 FILLER_1_2381 ();
 sg13g2_fill_1 FILLER_1_2385 ();
 sg13g2_decap_4 FILLER_1_2389 ();
 sg13g2_fill_1 FILLER_1_2393 ();
 sg13g2_decap_8 FILLER_1_2397 ();
 sg13g2_fill_2 FILLER_1_2404 ();
 sg13g2_decap_8 FILLER_1_2411 ();
 sg13g2_decap_8 FILLER_1_2418 ();
 sg13g2_decap_8 FILLER_1_2425 ();
 sg13g2_decap_4 FILLER_1_2432 ();
 sg13g2_fill_1 FILLER_1_2436 ();
 sg13g2_decap_8 FILLER_1_2442 ();
 sg13g2_decap_8 FILLER_1_2449 ();
 sg13g2_decap_8 FILLER_1_2456 ();
 sg13g2_decap_8 FILLER_1_2463 ();
 sg13g2_decap_8 FILLER_1_2470 ();
 sg13g2_decap_8 FILLER_1_2477 ();
 sg13g2_decap_8 FILLER_1_2484 ();
 sg13g2_decap_8 FILLER_1_2491 ();
 sg13g2_decap_8 FILLER_1_2498 ();
 sg13g2_decap_8 FILLER_1_2505 ();
 sg13g2_decap_4 FILLER_1_2512 ();
 sg13g2_fill_2 FILLER_1_2516 ();
 sg13g2_decap_8 FILLER_1_2523 ();
 sg13g2_decap_4 FILLER_1_2530 ();
 sg13g2_decap_4 FILLER_1_2540 ();
 sg13g2_fill_1 FILLER_1_2550 ();
 sg13g2_fill_2 FILLER_1_2557 ();
 sg13g2_fill_1 FILLER_1_2559 ();
 sg13g2_decap_4 FILLER_1_2572 ();
 sg13g2_fill_1 FILLER_1_2588 ();
 sg13g2_fill_2 FILLER_1_2595 ();
 sg13g2_fill_1 FILLER_1_2597 ();
 sg13g2_fill_2 FILLER_1_2610 ();
 sg13g2_fill_1 FILLER_1_2612 ();
 sg13g2_fill_2 FILLER_1_2619 ();
 sg13g2_fill_1 FILLER_1_2621 ();
 sg13g2_fill_2 FILLER_1_2634 ();
 sg13g2_fill_1 FILLER_1_2642 ();
 sg13g2_decap_4 FILLER_1_2649 ();
 sg13g2_fill_2 FILLER_1_2659 ();
 sg13g2_fill_1 FILLER_1_2661 ();
 sg13g2_decap_8 FILLER_1_2679 ();
 sg13g2_decap_8 FILLER_1_2686 ();
 sg13g2_decap_8 FILLER_1_2693 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_882 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_decap_8 FILLER_2_959 ();
 sg13g2_decap_8 FILLER_2_966 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_994 ();
 sg13g2_fill_2 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_2_1035 ();
 sg13g2_decap_4 FILLER_2_1042 ();
 sg13g2_fill_2 FILLER_2_1046 ();
 sg13g2_decap_8 FILLER_2_1073 ();
 sg13g2_decap_8 FILLER_2_1080 ();
 sg13g2_decap_4 FILLER_2_1087 ();
 sg13g2_fill_2 FILLER_2_1091 ();
 sg13g2_decap_8 FILLER_2_1114 ();
 sg13g2_decap_8 FILLER_2_1121 ();
 sg13g2_decap_8 FILLER_2_1128 ();
 sg13g2_decap_8 FILLER_2_1135 ();
 sg13g2_decap_8 FILLER_2_1142 ();
 sg13g2_decap_8 FILLER_2_1149 ();
 sg13g2_decap_8 FILLER_2_1156 ();
 sg13g2_decap_8 FILLER_2_1163 ();
 sg13g2_decap_8 FILLER_2_1170 ();
 sg13g2_decap_8 FILLER_2_1177 ();
 sg13g2_decap_8 FILLER_2_1184 ();
 sg13g2_decap_8 FILLER_2_1191 ();
 sg13g2_decap_8 FILLER_2_1198 ();
 sg13g2_decap_8 FILLER_2_1205 ();
 sg13g2_decap_8 FILLER_2_1212 ();
 sg13g2_decap_8 FILLER_2_1219 ();
 sg13g2_decap_8 FILLER_2_1226 ();
 sg13g2_decap_8 FILLER_2_1233 ();
 sg13g2_decap_8 FILLER_2_1240 ();
 sg13g2_decap_8 FILLER_2_1247 ();
 sg13g2_decap_8 FILLER_2_1254 ();
 sg13g2_decap_8 FILLER_2_1261 ();
 sg13g2_decap_8 FILLER_2_1268 ();
 sg13g2_decap_8 FILLER_2_1275 ();
 sg13g2_decap_8 FILLER_2_1282 ();
 sg13g2_decap_8 FILLER_2_1289 ();
 sg13g2_decap_8 FILLER_2_1296 ();
 sg13g2_decap_8 FILLER_2_1303 ();
 sg13g2_decap_8 FILLER_2_1310 ();
 sg13g2_decap_8 FILLER_2_1317 ();
 sg13g2_decap_8 FILLER_2_1324 ();
 sg13g2_decap_8 FILLER_2_1331 ();
 sg13g2_decap_8 FILLER_2_1338 ();
 sg13g2_decap_8 FILLER_2_1345 ();
 sg13g2_decap_8 FILLER_2_1352 ();
 sg13g2_decap_8 FILLER_2_1359 ();
 sg13g2_decap_8 FILLER_2_1366 ();
 sg13g2_decap_8 FILLER_2_1373 ();
 sg13g2_decap_8 FILLER_2_1380 ();
 sg13g2_decap_8 FILLER_2_1387 ();
 sg13g2_decap_8 FILLER_2_1394 ();
 sg13g2_decap_8 FILLER_2_1401 ();
 sg13g2_decap_8 FILLER_2_1408 ();
 sg13g2_decap_8 FILLER_2_1415 ();
 sg13g2_decap_8 FILLER_2_1422 ();
 sg13g2_decap_8 FILLER_2_1429 ();
 sg13g2_decap_8 FILLER_2_1436 ();
 sg13g2_decap_8 FILLER_2_1443 ();
 sg13g2_decap_8 FILLER_2_1450 ();
 sg13g2_decap_8 FILLER_2_1457 ();
 sg13g2_decap_8 FILLER_2_1464 ();
 sg13g2_decap_8 FILLER_2_1471 ();
 sg13g2_decap_8 FILLER_2_1478 ();
 sg13g2_decap_8 FILLER_2_1485 ();
 sg13g2_decap_8 FILLER_2_1492 ();
 sg13g2_decap_8 FILLER_2_1499 ();
 sg13g2_decap_8 FILLER_2_1506 ();
 sg13g2_decap_8 FILLER_2_1513 ();
 sg13g2_decap_8 FILLER_2_1520 ();
 sg13g2_decap_8 FILLER_2_1527 ();
 sg13g2_decap_8 FILLER_2_1534 ();
 sg13g2_decap_8 FILLER_2_1541 ();
 sg13g2_decap_8 FILLER_2_1548 ();
 sg13g2_decap_8 FILLER_2_1555 ();
 sg13g2_decap_8 FILLER_2_1562 ();
 sg13g2_decap_8 FILLER_2_1569 ();
 sg13g2_decap_8 FILLER_2_1576 ();
 sg13g2_decap_8 FILLER_2_1583 ();
 sg13g2_decap_8 FILLER_2_1590 ();
 sg13g2_decap_8 FILLER_2_1597 ();
 sg13g2_decap_8 FILLER_2_1604 ();
 sg13g2_decap_8 FILLER_2_1611 ();
 sg13g2_decap_8 FILLER_2_1618 ();
 sg13g2_decap_8 FILLER_2_1625 ();
 sg13g2_decap_8 FILLER_2_1632 ();
 sg13g2_decap_8 FILLER_2_1639 ();
 sg13g2_decap_8 FILLER_2_1646 ();
 sg13g2_decap_8 FILLER_2_1653 ();
 sg13g2_decap_8 FILLER_2_1660 ();
 sg13g2_decap_8 FILLER_2_1667 ();
 sg13g2_decap_8 FILLER_2_1674 ();
 sg13g2_decap_8 FILLER_2_1681 ();
 sg13g2_decap_8 FILLER_2_1688 ();
 sg13g2_decap_8 FILLER_2_1695 ();
 sg13g2_decap_8 FILLER_2_1702 ();
 sg13g2_decap_8 FILLER_2_1709 ();
 sg13g2_decap_8 FILLER_2_1716 ();
 sg13g2_decap_8 FILLER_2_1723 ();
 sg13g2_decap_8 FILLER_2_1730 ();
 sg13g2_decap_8 FILLER_2_1737 ();
 sg13g2_decap_8 FILLER_2_1744 ();
 sg13g2_decap_8 FILLER_2_1751 ();
 sg13g2_decap_8 FILLER_2_1758 ();
 sg13g2_decap_8 FILLER_2_1765 ();
 sg13g2_decap_8 FILLER_2_1772 ();
 sg13g2_decap_8 FILLER_2_1779 ();
 sg13g2_decap_8 FILLER_2_1786 ();
 sg13g2_decap_8 FILLER_2_1793 ();
 sg13g2_decap_8 FILLER_2_1800 ();
 sg13g2_decap_8 FILLER_2_1807 ();
 sg13g2_decap_8 FILLER_2_1814 ();
 sg13g2_decap_8 FILLER_2_1821 ();
 sg13g2_decap_8 FILLER_2_1828 ();
 sg13g2_decap_8 FILLER_2_1835 ();
 sg13g2_decap_8 FILLER_2_1842 ();
 sg13g2_decap_8 FILLER_2_1849 ();
 sg13g2_decap_8 FILLER_2_1856 ();
 sg13g2_decap_8 FILLER_2_1863 ();
 sg13g2_decap_8 FILLER_2_1870 ();
 sg13g2_decap_8 FILLER_2_1877 ();
 sg13g2_decap_8 FILLER_2_1884 ();
 sg13g2_decap_8 FILLER_2_1891 ();
 sg13g2_decap_4 FILLER_2_1898 ();
 sg13g2_fill_2 FILLER_2_1902 ();
 sg13g2_decap_8 FILLER_2_1929 ();
 sg13g2_decap_8 FILLER_2_1936 ();
 sg13g2_decap_4 FILLER_2_1943 ();
 sg13g2_decap_8 FILLER_2_1968 ();
 sg13g2_decap_8 FILLER_2_1975 ();
 sg13g2_decap_4 FILLER_2_1982 ();
 sg13g2_decap_8 FILLER_2_2007 ();
 sg13g2_decap_8 FILLER_2_2014 ();
 sg13g2_decap_8 FILLER_2_2021 ();
 sg13g2_fill_1 FILLER_2_2028 ();
 sg13g2_decap_8 FILLER_2_2050 ();
 sg13g2_decap_8 FILLER_2_2057 ();
 sg13g2_decap_8 FILLER_2_2064 ();
 sg13g2_decap_8 FILLER_2_2071 ();
 sg13g2_decap_8 FILLER_2_2078 ();
 sg13g2_decap_8 FILLER_2_2085 ();
 sg13g2_decap_8 FILLER_2_2092 ();
 sg13g2_fill_2 FILLER_2_2099 ();
 sg13g2_fill_1 FILLER_2_2101 ();
 sg13g2_decap_8 FILLER_2_2105 ();
 sg13g2_decap_8 FILLER_2_2112 ();
 sg13g2_decap_8 FILLER_2_2119 ();
 sg13g2_decap_8 FILLER_2_2126 ();
 sg13g2_decap_8 FILLER_2_2133 ();
 sg13g2_decap_8 FILLER_2_2140 ();
 sg13g2_fill_1 FILLER_2_2147 ();
 sg13g2_decap_8 FILLER_2_2151 ();
 sg13g2_decap_8 FILLER_2_2158 ();
 sg13g2_decap_8 FILLER_2_2165 ();
 sg13g2_decap_8 FILLER_2_2172 ();
 sg13g2_decap_4 FILLER_2_2179 ();
 sg13g2_fill_2 FILLER_2_2183 ();
 sg13g2_decap_8 FILLER_2_2188 ();
 sg13g2_decap_8 FILLER_2_2195 ();
 sg13g2_decap_8 FILLER_2_2202 ();
 sg13g2_decap_8 FILLER_2_2209 ();
 sg13g2_decap_8 FILLER_2_2219 ();
 sg13g2_decap_8 FILLER_2_2226 ();
 sg13g2_decap_8 FILLER_2_2233 ();
 sg13g2_decap_8 FILLER_2_2240 ();
 sg13g2_decap_8 FILLER_2_2247 ();
 sg13g2_decap_8 FILLER_2_2254 ();
 sg13g2_decap_8 FILLER_2_2261 ();
 sg13g2_fill_2 FILLER_2_2268 ();
 sg13g2_decap_8 FILLER_2_2285 ();
 sg13g2_decap_4 FILLER_2_2292 ();
 sg13g2_fill_1 FILLER_2_2296 ();
 sg13g2_decap_8 FILLER_2_2342 ();
 sg13g2_decap_4 FILLER_2_2349 ();
 sg13g2_fill_1 FILLER_2_2353 ();
 sg13g2_decap_8 FILLER_2_2379 ();
 sg13g2_decap_8 FILLER_2_2386 ();
 sg13g2_fill_2 FILLER_2_2393 ();
 sg13g2_fill_1 FILLER_2_2395 ();
 sg13g2_decap_4 FILLER_2_2421 ();
 sg13g2_fill_2 FILLER_2_2425 ();
 sg13g2_decap_4 FILLER_2_2502 ();
 sg13g2_fill_1 FILLER_2_2506 ();
 sg13g2_decap_8 FILLER_2_2532 ();
 sg13g2_decap_8 FILLER_2_2539 ();
 sg13g2_decap_8 FILLER_2_2546 ();
 sg13g2_decap_8 FILLER_2_2553 ();
 sg13g2_decap_8 FILLER_2_2560 ();
 sg13g2_decap_8 FILLER_2_2567 ();
 sg13g2_decap_8 FILLER_2_2574 ();
 sg13g2_decap_8 FILLER_2_2581 ();
 sg13g2_decap_8 FILLER_2_2588 ();
 sg13g2_decap_8 FILLER_2_2595 ();
 sg13g2_decap_8 FILLER_2_2602 ();
 sg13g2_decap_8 FILLER_2_2609 ();
 sg13g2_decap_8 FILLER_2_2616 ();
 sg13g2_decap_8 FILLER_2_2623 ();
 sg13g2_decap_8 FILLER_2_2630 ();
 sg13g2_decap_8 FILLER_2_2637 ();
 sg13g2_decap_8 FILLER_2_2644 ();
 sg13g2_decap_8 FILLER_2_2651 ();
 sg13g2_decap_8 FILLER_2_2658 ();
 sg13g2_decap_8 FILLER_2_2665 ();
 sg13g2_decap_8 FILLER_2_2672 ();
 sg13g2_decap_4 FILLER_2_2679 ();
 sg13g2_decap_8 FILLER_2_2687 ();
 sg13g2_decap_4 FILLER_2_2694 ();
 sg13g2_fill_2 FILLER_2_2698 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_fill_2 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_548 ();
 sg13g2_decap_8 FILLER_3_555 ();
 sg13g2_decap_8 FILLER_3_562 ();
 sg13g2_decap_8 FILLER_3_569 ();
 sg13g2_decap_8 FILLER_3_576 ();
 sg13g2_decap_8 FILLER_3_583 ();
 sg13g2_decap_8 FILLER_3_590 ();
 sg13g2_decap_8 FILLER_3_597 ();
 sg13g2_decap_8 FILLER_3_604 ();
 sg13g2_decap_8 FILLER_3_611 ();
 sg13g2_decap_8 FILLER_3_618 ();
 sg13g2_decap_8 FILLER_3_625 ();
 sg13g2_decap_8 FILLER_3_632 ();
 sg13g2_decap_8 FILLER_3_639 ();
 sg13g2_decap_8 FILLER_3_646 ();
 sg13g2_decap_8 FILLER_3_653 ();
 sg13g2_decap_8 FILLER_3_660 ();
 sg13g2_decap_8 FILLER_3_667 ();
 sg13g2_decap_8 FILLER_3_674 ();
 sg13g2_decap_8 FILLER_3_681 ();
 sg13g2_decap_8 FILLER_3_688 ();
 sg13g2_decap_8 FILLER_3_695 ();
 sg13g2_decap_8 FILLER_3_702 ();
 sg13g2_decap_8 FILLER_3_709 ();
 sg13g2_decap_8 FILLER_3_716 ();
 sg13g2_decap_8 FILLER_3_723 ();
 sg13g2_decap_8 FILLER_3_730 ();
 sg13g2_decap_8 FILLER_3_737 ();
 sg13g2_decap_8 FILLER_3_744 ();
 sg13g2_decap_8 FILLER_3_751 ();
 sg13g2_decap_8 FILLER_3_758 ();
 sg13g2_decap_8 FILLER_3_765 ();
 sg13g2_decap_8 FILLER_3_772 ();
 sg13g2_decap_8 FILLER_3_779 ();
 sg13g2_decap_8 FILLER_3_786 ();
 sg13g2_decap_8 FILLER_3_793 ();
 sg13g2_fill_2 FILLER_3_800 ();
 sg13g2_decap_8 FILLER_3_827 ();
 sg13g2_decap_8 FILLER_3_834 ();
 sg13g2_fill_2 FILLER_3_841 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_decap_8 FILLER_3_875 ();
 sg13g2_decap_8 FILLER_3_882 ();
 sg13g2_decap_8 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_910 ();
 sg13g2_decap_8 FILLER_3_917 ();
 sg13g2_decap_8 FILLER_3_924 ();
 sg13g2_decap_8 FILLER_3_931 ();
 sg13g2_decap_8 FILLER_3_938 ();
 sg13g2_decap_8 FILLER_3_945 ();
 sg13g2_decap_8 FILLER_3_952 ();
 sg13g2_decap_8 FILLER_3_959 ();
 sg13g2_decap_4 FILLER_3_966 ();
 sg13g2_decap_8 FILLER_3_983 ();
 sg13g2_decap_8 FILLER_3_990 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_8 FILLER_3_1025 ();
 sg13g2_decap_8 FILLER_3_1032 ();
 sg13g2_decap_8 FILLER_3_1039 ();
 sg13g2_decap_8 FILLER_3_1046 ();
 sg13g2_decap_8 FILLER_3_1053 ();
 sg13g2_decap_8 FILLER_3_1060 ();
 sg13g2_decap_8 FILLER_3_1067 ();
 sg13g2_decap_8 FILLER_3_1074 ();
 sg13g2_decap_8 FILLER_3_1081 ();
 sg13g2_fill_2 FILLER_3_1088 ();
 sg13g2_decap_8 FILLER_3_1115 ();
 sg13g2_decap_8 FILLER_3_1122 ();
 sg13g2_decap_4 FILLER_3_1129 ();
 sg13g2_decap_8 FILLER_3_1154 ();
 sg13g2_decap_8 FILLER_3_1161 ();
 sg13g2_decap_4 FILLER_3_1168 ();
 sg13g2_fill_1 FILLER_3_1172 ();
 sg13g2_decap_8 FILLER_3_1194 ();
 sg13g2_decap_8 FILLER_3_1201 ();
 sg13g2_decap_8 FILLER_3_1208 ();
 sg13g2_fill_2 FILLER_3_1215 ();
 sg13g2_decap_8 FILLER_3_1220 ();
 sg13g2_decap_8 FILLER_3_1227 ();
 sg13g2_decap_8 FILLER_3_1234 ();
 sg13g2_decap_8 FILLER_3_1241 ();
 sg13g2_decap_8 FILLER_3_1248 ();
 sg13g2_decap_8 FILLER_3_1255 ();
 sg13g2_decap_8 FILLER_3_1262 ();
 sg13g2_decap_8 FILLER_3_1269 ();
 sg13g2_decap_8 FILLER_3_1276 ();
 sg13g2_decap_8 FILLER_3_1283 ();
 sg13g2_decap_8 FILLER_3_1290 ();
 sg13g2_decap_8 FILLER_3_1297 ();
 sg13g2_decap_8 FILLER_3_1304 ();
 sg13g2_decap_8 FILLER_3_1311 ();
 sg13g2_decap_8 FILLER_3_1318 ();
 sg13g2_decap_8 FILLER_3_1325 ();
 sg13g2_fill_2 FILLER_3_1332 ();
 sg13g2_decap_8 FILLER_3_1347 ();
 sg13g2_decap_8 FILLER_3_1354 ();
 sg13g2_decap_8 FILLER_3_1361 ();
 sg13g2_decap_8 FILLER_3_1368 ();
 sg13g2_decap_8 FILLER_3_1375 ();
 sg13g2_decap_8 FILLER_3_1382 ();
 sg13g2_decap_8 FILLER_3_1389 ();
 sg13g2_decap_8 FILLER_3_1396 ();
 sg13g2_decap_8 FILLER_3_1403 ();
 sg13g2_decap_8 FILLER_3_1410 ();
 sg13g2_decap_8 FILLER_3_1417 ();
 sg13g2_decap_8 FILLER_3_1424 ();
 sg13g2_decap_4 FILLER_3_1431 ();
 sg13g2_fill_2 FILLER_3_1435 ();
 sg13g2_decap_8 FILLER_3_1440 ();
 sg13g2_decap_8 FILLER_3_1447 ();
 sg13g2_decap_8 FILLER_3_1454 ();
 sg13g2_decap_8 FILLER_3_1461 ();
 sg13g2_decap_8 FILLER_3_1468 ();
 sg13g2_decap_8 FILLER_3_1475 ();
 sg13g2_decap_8 FILLER_3_1482 ();
 sg13g2_decap_8 FILLER_3_1489 ();
 sg13g2_decap_8 FILLER_3_1496 ();
 sg13g2_decap_8 FILLER_3_1503 ();
 sg13g2_decap_8 FILLER_3_1510 ();
 sg13g2_decap_8 FILLER_3_1517 ();
 sg13g2_decap_8 FILLER_3_1524 ();
 sg13g2_decap_8 FILLER_3_1531 ();
 sg13g2_decap_8 FILLER_3_1538 ();
 sg13g2_decap_8 FILLER_3_1545 ();
 sg13g2_decap_8 FILLER_3_1552 ();
 sg13g2_decap_8 FILLER_3_1559 ();
 sg13g2_decap_8 FILLER_3_1566 ();
 sg13g2_decap_8 FILLER_3_1573 ();
 sg13g2_decap_8 FILLER_3_1580 ();
 sg13g2_decap_8 FILLER_3_1587 ();
 sg13g2_decap_8 FILLER_3_1594 ();
 sg13g2_decap_8 FILLER_3_1601 ();
 sg13g2_decap_8 FILLER_3_1608 ();
 sg13g2_decap_8 FILLER_3_1615 ();
 sg13g2_decap_8 FILLER_3_1622 ();
 sg13g2_decap_8 FILLER_3_1629 ();
 sg13g2_decap_8 FILLER_3_1636 ();
 sg13g2_decap_8 FILLER_3_1643 ();
 sg13g2_decap_8 FILLER_3_1650 ();
 sg13g2_decap_8 FILLER_3_1657 ();
 sg13g2_decap_8 FILLER_3_1664 ();
 sg13g2_decap_8 FILLER_3_1671 ();
 sg13g2_decap_8 FILLER_3_1678 ();
 sg13g2_decap_8 FILLER_3_1685 ();
 sg13g2_decap_8 FILLER_3_1692 ();
 sg13g2_decap_8 FILLER_3_1699 ();
 sg13g2_decap_8 FILLER_3_1706 ();
 sg13g2_decap_8 FILLER_3_1713 ();
 sg13g2_decap_8 FILLER_3_1720 ();
 sg13g2_decap_8 FILLER_3_1727 ();
 sg13g2_decap_8 FILLER_3_1734 ();
 sg13g2_decap_8 FILLER_3_1741 ();
 sg13g2_decap_8 FILLER_3_1761 ();
 sg13g2_decap_8 FILLER_3_1768 ();
 sg13g2_decap_8 FILLER_3_1775 ();
 sg13g2_decap_8 FILLER_3_1782 ();
 sg13g2_decap_8 FILLER_3_1789 ();
 sg13g2_decap_4 FILLER_3_1796 ();
 sg13g2_fill_2 FILLER_3_1800 ();
 sg13g2_decap_8 FILLER_3_1815 ();
 sg13g2_decap_8 FILLER_3_1822 ();
 sg13g2_decap_8 FILLER_3_1829 ();
 sg13g2_decap_8 FILLER_3_1836 ();
 sg13g2_decap_8 FILLER_3_1843 ();
 sg13g2_decap_8 FILLER_3_1850 ();
 sg13g2_decap_8 FILLER_3_1857 ();
 sg13g2_decap_8 FILLER_3_1864 ();
 sg13g2_decap_8 FILLER_3_1871 ();
 sg13g2_decap_8 FILLER_3_1878 ();
 sg13g2_decap_8 FILLER_3_1885 ();
 sg13g2_decap_8 FILLER_3_1892 ();
 sg13g2_decap_8 FILLER_3_1899 ();
 sg13g2_decap_8 FILLER_3_1906 ();
 sg13g2_decap_8 FILLER_3_1913 ();
 sg13g2_decap_8 FILLER_3_1920 ();
 sg13g2_decap_8 FILLER_3_1927 ();
 sg13g2_decap_8 FILLER_3_1934 ();
 sg13g2_fill_2 FILLER_3_1941 ();
 sg13g2_fill_1 FILLER_3_1943 ();
 sg13g2_decap_8 FILLER_3_1969 ();
 sg13g2_decap_8 FILLER_3_1976 ();
 sg13g2_fill_1 FILLER_3_1983 ();
 sg13g2_decap_8 FILLER_3_2009 ();
 sg13g2_decap_8 FILLER_3_2016 ();
 sg13g2_fill_1 FILLER_3_2023 ();
 sg13g2_decap_8 FILLER_3_2049 ();
 sg13g2_decap_8 FILLER_3_2056 ();
 sg13g2_decap_8 FILLER_3_2084 ();
 sg13g2_decap_8 FILLER_3_2091 ();
 sg13g2_decap_8 FILLER_3_2098 ();
 sg13g2_decap_8 FILLER_3_2105 ();
 sg13g2_decap_8 FILLER_3_2112 ();
 sg13g2_decap_8 FILLER_3_2119 ();
 sg13g2_decap_8 FILLER_3_2126 ();
 sg13g2_fill_1 FILLER_3_2133 ();
 sg13g2_fill_2 FILLER_3_2137 ();
 sg13g2_fill_1 FILLER_3_2139 ();
 sg13g2_decap_8 FILLER_3_2143 ();
 sg13g2_decap_8 FILLER_3_2150 ();
 sg13g2_decap_8 FILLER_3_2157 ();
 sg13g2_decap_8 FILLER_3_2164 ();
 sg13g2_decap_8 FILLER_3_2171 ();
 sg13g2_decap_8 FILLER_3_2178 ();
 sg13g2_decap_8 FILLER_3_2185 ();
 sg13g2_decap_8 FILLER_3_2192 ();
 sg13g2_decap_8 FILLER_3_2199 ();
 sg13g2_decap_8 FILLER_3_2206 ();
 sg13g2_decap_8 FILLER_3_2213 ();
 sg13g2_decap_8 FILLER_3_2220 ();
 sg13g2_decap_8 FILLER_3_2227 ();
 sg13g2_decap_8 FILLER_3_2234 ();
 sg13g2_fill_2 FILLER_3_2241 ();
 sg13g2_fill_1 FILLER_3_2243 ();
 sg13g2_decap_8 FILLER_3_2257 ();
 sg13g2_decap_8 FILLER_3_2264 ();
 sg13g2_decap_8 FILLER_3_2271 ();
 sg13g2_decap_8 FILLER_3_2278 ();
 sg13g2_decap_8 FILLER_3_2285 ();
 sg13g2_decap_8 FILLER_3_2292 ();
 sg13g2_decap_8 FILLER_3_2299 ();
 sg13g2_decap_8 FILLER_3_2306 ();
 sg13g2_decap_8 FILLER_3_2313 ();
 sg13g2_decap_8 FILLER_3_2320 ();
 sg13g2_decap_8 FILLER_3_2327 ();
 sg13g2_decap_8 FILLER_3_2334 ();
 sg13g2_decap_8 FILLER_3_2341 ();
 sg13g2_decap_8 FILLER_3_2348 ();
 sg13g2_decap_8 FILLER_3_2355 ();
 sg13g2_decap_8 FILLER_3_2362 ();
 sg13g2_decap_8 FILLER_3_2369 ();
 sg13g2_decap_8 FILLER_3_2376 ();
 sg13g2_decap_8 FILLER_3_2383 ();
 sg13g2_decap_8 FILLER_3_2390 ();
 sg13g2_decap_8 FILLER_3_2397 ();
 sg13g2_decap_8 FILLER_3_2404 ();
 sg13g2_decap_8 FILLER_3_2411 ();
 sg13g2_decap_8 FILLER_3_2418 ();
 sg13g2_decap_8 FILLER_3_2425 ();
 sg13g2_decap_8 FILLER_3_2432 ();
 sg13g2_decap_8 FILLER_3_2439 ();
 sg13g2_decap_8 FILLER_3_2446 ();
 sg13g2_decap_8 FILLER_3_2453 ();
 sg13g2_decap_8 FILLER_3_2460 ();
 sg13g2_decap_8 FILLER_3_2467 ();
 sg13g2_decap_8 FILLER_3_2474 ();
 sg13g2_fill_2 FILLER_3_2481 ();
 sg13g2_fill_1 FILLER_3_2483 ();
 sg13g2_decap_8 FILLER_3_2489 ();
 sg13g2_decap_8 FILLER_3_2496 ();
 sg13g2_decap_8 FILLER_3_2503 ();
 sg13g2_decap_8 FILLER_3_2510 ();
 sg13g2_decap_8 FILLER_3_2517 ();
 sg13g2_decap_8 FILLER_3_2524 ();
 sg13g2_decap_8 FILLER_3_2531 ();
 sg13g2_decap_8 FILLER_3_2538 ();
 sg13g2_decap_8 FILLER_3_2545 ();
 sg13g2_decap_8 FILLER_3_2552 ();
 sg13g2_decap_8 FILLER_3_2559 ();
 sg13g2_decap_8 FILLER_3_2566 ();
 sg13g2_decap_8 FILLER_3_2573 ();
 sg13g2_decap_8 FILLER_3_2580 ();
 sg13g2_decap_8 FILLER_3_2587 ();
 sg13g2_decap_8 FILLER_3_2594 ();
 sg13g2_decap_8 FILLER_3_2601 ();
 sg13g2_decap_8 FILLER_3_2608 ();
 sg13g2_decap_8 FILLER_3_2615 ();
 sg13g2_decap_8 FILLER_3_2622 ();
 sg13g2_decap_8 FILLER_3_2629 ();
 sg13g2_decap_8 FILLER_3_2636 ();
 sg13g2_decap_8 FILLER_3_2643 ();
 sg13g2_decap_8 FILLER_3_2650 ();
 sg13g2_decap_8 FILLER_3_2657 ();
 sg13g2_decap_8 FILLER_3_2664 ();
 sg13g2_decap_8 FILLER_3_2671 ();
 sg13g2_decap_8 FILLER_3_2678 ();
 sg13g2_decap_8 FILLER_3_2685 ();
 sg13g2_decap_8 FILLER_3_2692 ();
 sg13g2_fill_1 FILLER_3_2699 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_fill_1 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_554 ();
 sg13g2_decap_8 FILLER_4_561 ();
 sg13g2_decap_4 FILLER_4_568 ();
 sg13g2_fill_1 FILLER_4_572 ();
 sg13g2_decap_8 FILLER_4_615 ();
 sg13g2_decap_8 FILLER_4_622 ();
 sg13g2_decap_8 FILLER_4_629 ();
 sg13g2_decap_8 FILLER_4_636 ();
 sg13g2_decap_8 FILLER_4_643 ();
 sg13g2_decap_8 FILLER_4_650 ();
 sg13g2_decap_8 FILLER_4_657 ();
 sg13g2_decap_4 FILLER_4_664 ();
 sg13g2_decap_8 FILLER_4_689 ();
 sg13g2_decap_8 FILLER_4_696 ();
 sg13g2_decap_8 FILLER_4_703 ();
 sg13g2_decap_8 FILLER_4_710 ();
 sg13g2_decap_8 FILLER_4_717 ();
 sg13g2_decap_8 FILLER_4_724 ();
 sg13g2_decap_8 FILLER_4_731 ();
 sg13g2_fill_2 FILLER_4_738 ();
 sg13g2_decap_8 FILLER_4_765 ();
 sg13g2_decap_8 FILLER_4_772 ();
 sg13g2_decap_8 FILLER_4_779 ();
 sg13g2_decap_8 FILLER_4_786 ();
 sg13g2_decap_8 FILLER_4_793 ();
 sg13g2_decap_8 FILLER_4_800 ();
 sg13g2_decap_8 FILLER_4_807 ();
 sg13g2_decap_8 FILLER_4_814 ();
 sg13g2_decap_8 FILLER_4_821 ();
 sg13g2_decap_8 FILLER_4_828 ();
 sg13g2_decap_8 FILLER_4_835 ();
 sg13g2_decap_8 FILLER_4_842 ();
 sg13g2_decap_8 FILLER_4_849 ();
 sg13g2_decap_8 FILLER_4_856 ();
 sg13g2_decap_8 FILLER_4_863 ();
 sg13g2_decap_4 FILLER_4_870 ();
 sg13g2_fill_2 FILLER_4_874 ();
 sg13g2_decap_4 FILLER_4_889 ();
 sg13g2_fill_2 FILLER_4_893 ();
 sg13g2_decap_8 FILLER_4_920 ();
 sg13g2_decap_4 FILLER_4_927 ();
 sg13g2_fill_1 FILLER_4_931 ();
 sg13g2_decap_8 FILLER_4_957 ();
 sg13g2_decap_8 FILLER_4_964 ();
 sg13g2_fill_2 FILLER_4_971 ();
 sg13g2_fill_1 FILLER_4_973 ();
 sg13g2_decap_8 FILLER_4_984 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_8 FILLER_4_1005 ();
 sg13g2_decap_8 FILLER_4_1012 ();
 sg13g2_decap_8 FILLER_4_1019 ();
 sg13g2_decap_8 FILLER_4_1026 ();
 sg13g2_decap_8 FILLER_4_1033 ();
 sg13g2_decap_8 FILLER_4_1040 ();
 sg13g2_decap_8 FILLER_4_1047 ();
 sg13g2_decap_8 FILLER_4_1054 ();
 sg13g2_decap_8 FILLER_4_1061 ();
 sg13g2_decap_8 FILLER_4_1068 ();
 sg13g2_decap_8 FILLER_4_1075 ();
 sg13g2_decap_8 FILLER_4_1082 ();
 sg13g2_decap_8 FILLER_4_1089 ();
 sg13g2_decap_8 FILLER_4_1096 ();
 sg13g2_decap_8 FILLER_4_1103 ();
 sg13g2_decap_8 FILLER_4_1110 ();
 sg13g2_decap_8 FILLER_4_1117 ();
 sg13g2_decap_8 FILLER_4_1124 ();
 sg13g2_decap_8 FILLER_4_1156 ();
 sg13g2_decap_8 FILLER_4_1163 ();
 sg13g2_fill_1 FILLER_4_1170 ();
 sg13g2_decap_8 FILLER_4_1196 ();
 sg13g2_decap_8 FILLER_4_1203 ();
 sg13g2_decap_8 FILLER_4_1210 ();
 sg13g2_decap_8 FILLER_4_1217 ();
 sg13g2_decap_8 FILLER_4_1224 ();
 sg13g2_decap_8 FILLER_4_1231 ();
 sg13g2_decap_8 FILLER_4_1238 ();
 sg13g2_decap_8 FILLER_4_1245 ();
 sg13g2_decap_4 FILLER_4_1252 ();
 sg13g2_decap_8 FILLER_4_1277 ();
 sg13g2_decap_8 FILLER_4_1284 ();
 sg13g2_decap_8 FILLER_4_1291 ();
 sg13g2_fill_2 FILLER_4_1298 ();
 sg13g2_fill_1 FILLER_4_1300 ();
 sg13g2_decap_8 FILLER_4_1322 ();
 sg13g2_decap_4 FILLER_4_1329 ();
 sg13g2_fill_2 FILLER_4_1333 ();
 sg13g2_decap_8 FILLER_4_1340 ();
 sg13g2_decap_8 FILLER_4_1347 ();
 sg13g2_decap_8 FILLER_4_1354 ();
 sg13g2_decap_8 FILLER_4_1361 ();
 sg13g2_decap_8 FILLER_4_1368 ();
 sg13g2_decap_8 FILLER_4_1375 ();
 sg13g2_decap_8 FILLER_4_1382 ();
 sg13g2_decap_8 FILLER_4_1389 ();
 sg13g2_decap_8 FILLER_4_1396 ();
 sg13g2_decap_8 FILLER_4_1403 ();
 sg13g2_decap_8 FILLER_4_1410 ();
 sg13g2_decap_8 FILLER_4_1417 ();
 sg13g2_decap_8 FILLER_4_1424 ();
 sg13g2_decap_8 FILLER_4_1431 ();
 sg13g2_decap_8 FILLER_4_1438 ();
 sg13g2_decap_8 FILLER_4_1445 ();
 sg13g2_decap_8 FILLER_4_1452 ();
 sg13g2_decap_8 FILLER_4_1459 ();
 sg13g2_decap_8 FILLER_4_1466 ();
 sg13g2_decap_4 FILLER_4_1473 ();
 sg13g2_fill_1 FILLER_4_1477 ();
 sg13g2_decap_8 FILLER_4_1481 ();
 sg13g2_decap_8 FILLER_4_1488 ();
 sg13g2_decap_8 FILLER_4_1495 ();
 sg13g2_decap_8 FILLER_4_1502 ();
 sg13g2_decap_8 FILLER_4_1509 ();
 sg13g2_decap_8 FILLER_4_1516 ();
 sg13g2_decap_8 FILLER_4_1523 ();
 sg13g2_decap_8 FILLER_4_1530 ();
 sg13g2_decap_8 FILLER_4_1537 ();
 sg13g2_decap_8 FILLER_4_1544 ();
 sg13g2_decap_8 FILLER_4_1551 ();
 sg13g2_decap_8 FILLER_4_1558 ();
 sg13g2_decap_8 FILLER_4_1565 ();
 sg13g2_decap_8 FILLER_4_1572 ();
 sg13g2_decap_8 FILLER_4_1579 ();
 sg13g2_decap_8 FILLER_4_1586 ();
 sg13g2_decap_8 FILLER_4_1593 ();
 sg13g2_decap_8 FILLER_4_1600 ();
 sg13g2_decap_8 FILLER_4_1607 ();
 sg13g2_decap_8 FILLER_4_1614 ();
 sg13g2_decap_8 FILLER_4_1621 ();
 sg13g2_decap_8 FILLER_4_1628 ();
 sg13g2_decap_8 FILLER_4_1635 ();
 sg13g2_decap_8 FILLER_4_1642 ();
 sg13g2_decap_8 FILLER_4_1649 ();
 sg13g2_decap_8 FILLER_4_1656 ();
 sg13g2_decap_8 FILLER_4_1663 ();
 sg13g2_decap_8 FILLER_4_1670 ();
 sg13g2_decap_8 FILLER_4_1677 ();
 sg13g2_decap_8 FILLER_4_1684 ();
 sg13g2_decap_8 FILLER_4_1691 ();
 sg13g2_decap_8 FILLER_4_1698 ();
 sg13g2_decap_8 FILLER_4_1705 ();
 sg13g2_decap_8 FILLER_4_1712 ();
 sg13g2_decap_8 FILLER_4_1719 ();
 sg13g2_decap_8 FILLER_4_1726 ();
 sg13g2_decap_8 FILLER_4_1733 ();
 sg13g2_decap_4 FILLER_4_1740 ();
 sg13g2_fill_2 FILLER_4_1744 ();
 sg13g2_decap_8 FILLER_4_1751 ();
 sg13g2_decap_8 FILLER_4_1758 ();
 sg13g2_decap_8 FILLER_4_1765 ();
 sg13g2_decap_8 FILLER_4_1772 ();
 sg13g2_decap_8 FILLER_4_1779 ();
 sg13g2_decap_8 FILLER_4_1786 ();
 sg13g2_fill_2 FILLER_4_1793 ();
 sg13g2_fill_1 FILLER_4_1795 ();
 sg13g2_decap_8 FILLER_4_1801 ();
 sg13g2_decap_8 FILLER_4_1808 ();
 sg13g2_decap_8 FILLER_4_1815 ();
 sg13g2_decap_8 FILLER_4_1822 ();
 sg13g2_decap_8 FILLER_4_1829 ();
 sg13g2_decap_8 FILLER_4_1836 ();
 sg13g2_decap_8 FILLER_4_1843 ();
 sg13g2_decap_8 FILLER_4_1850 ();
 sg13g2_decap_8 FILLER_4_1857 ();
 sg13g2_decap_8 FILLER_4_1864 ();
 sg13g2_decap_8 FILLER_4_1871 ();
 sg13g2_decap_8 FILLER_4_1878 ();
 sg13g2_decap_8 FILLER_4_1885 ();
 sg13g2_decap_8 FILLER_4_1892 ();
 sg13g2_decap_8 FILLER_4_1899 ();
 sg13g2_decap_8 FILLER_4_1906 ();
 sg13g2_decap_8 FILLER_4_1913 ();
 sg13g2_decap_8 FILLER_4_1920 ();
 sg13g2_decap_8 FILLER_4_1927 ();
 sg13g2_decap_8 FILLER_4_1934 ();
 sg13g2_decap_8 FILLER_4_1941 ();
 sg13g2_decap_8 FILLER_4_1948 ();
 sg13g2_decap_8 FILLER_4_1955 ();
 sg13g2_decap_8 FILLER_4_1962 ();
 sg13g2_decap_8 FILLER_4_1969 ();
 sg13g2_decap_8 FILLER_4_1976 ();
 sg13g2_decap_8 FILLER_4_1983 ();
 sg13g2_decap_8 FILLER_4_1990 ();
 sg13g2_decap_8 FILLER_4_1997 ();
 sg13g2_decap_8 FILLER_4_2004 ();
 sg13g2_decap_8 FILLER_4_2011 ();
 sg13g2_decap_8 FILLER_4_2018 ();
 sg13g2_decap_8 FILLER_4_2025 ();
 sg13g2_decap_8 FILLER_4_2032 ();
 sg13g2_decap_8 FILLER_4_2039 ();
 sg13g2_decap_8 FILLER_4_2046 ();
 sg13g2_decap_8 FILLER_4_2053 ();
 sg13g2_fill_1 FILLER_4_2060 ();
 sg13g2_decap_8 FILLER_4_2086 ();
 sg13g2_decap_8 FILLER_4_2093 ();
 sg13g2_decap_8 FILLER_4_2100 ();
 sg13g2_decap_4 FILLER_4_2107 ();
 sg13g2_fill_2 FILLER_4_2111 ();
 sg13g2_decap_8 FILLER_4_2116 ();
 sg13g2_decap_8 FILLER_4_2123 ();
 sg13g2_decap_8 FILLER_4_2130 ();
 sg13g2_decap_8 FILLER_4_2137 ();
 sg13g2_decap_8 FILLER_4_2144 ();
 sg13g2_decap_8 FILLER_4_2151 ();
 sg13g2_decap_8 FILLER_4_2158 ();
 sg13g2_decap_4 FILLER_4_2165 ();
 sg13g2_fill_1 FILLER_4_2169 ();
 sg13g2_decap_8 FILLER_4_2191 ();
 sg13g2_decap_8 FILLER_4_2198 ();
 sg13g2_decap_4 FILLER_4_2205 ();
 sg13g2_fill_2 FILLER_4_2209 ();
 sg13g2_fill_2 FILLER_4_2232 ();
 sg13g2_fill_1 FILLER_4_2234 ();
 sg13g2_decap_8 FILLER_4_2240 ();
 sg13g2_decap_8 FILLER_4_2247 ();
 sg13g2_decap_8 FILLER_4_2254 ();
 sg13g2_decap_8 FILLER_4_2261 ();
 sg13g2_decap_8 FILLER_4_2268 ();
 sg13g2_decap_8 FILLER_4_2275 ();
 sg13g2_decap_8 FILLER_4_2282 ();
 sg13g2_decap_8 FILLER_4_2289 ();
 sg13g2_decap_8 FILLER_4_2296 ();
 sg13g2_decap_8 FILLER_4_2303 ();
 sg13g2_decap_8 FILLER_4_2310 ();
 sg13g2_decap_8 FILLER_4_2317 ();
 sg13g2_decap_8 FILLER_4_2324 ();
 sg13g2_decap_8 FILLER_4_2331 ();
 sg13g2_decap_8 FILLER_4_2338 ();
 sg13g2_decap_8 FILLER_4_2345 ();
 sg13g2_decap_8 FILLER_4_2352 ();
 sg13g2_decap_8 FILLER_4_2364 ();
 sg13g2_decap_8 FILLER_4_2371 ();
 sg13g2_decap_8 FILLER_4_2378 ();
 sg13g2_decap_8 FILLER_4_2385 ();
 sg13g2_decap_8 FILLER_4_2392 ();
 sg13g2_decap_8 FILLER_4_2399 ();
 sg13g2_decap_8 FILLER_4_2406 ();
 sg13g2_decap_8 FILLER_4_2413 ();
 sg13g2_decap_8 FILLER_4_2420 ();
 sg13g2_fill_2 FILLER_4_2427 ();
 sg13g2_decap_8 FILLER_4_2434 ();
 sg13g2_decap_8 FILLER_4_2441 ();
 sg13g2_decap_8 FILLER_4_2448 ();
 sg13g2_decap_8 FILLER_4_2455 ();
 sg13g2_fill_1 FILLER_4_2462 ();
 sg13g2_decap_8 FILLER_4_2468 ();
 sg13g2_decap_8 FILLER_4_2475 ();
 sg13g2_decap_8 FILLER_4_2482 ();
 sg13g2_decap_8 FILLER_4_2489 ();
 sg13g2_decap_8 FILLER_4_2496 ();
 sg13g2_decap_8 FILLER_4_2503 ();
 sg13g2_decap_8 FILLER_4_2510 ();
 sg13g2_decap_8 FILLER_4_2517 ();
 sg13g2_fill_2 FILLER_4_2524 ();
 sg13g2_decap_8 FILLER_4_2551 ();
 sg13g2_decap_8 FILLER_4_2558 ();
 sg13g2_decap_8 FILLER_4_2565 ();
 sg13g2_decap_8 FILLER_4_2572 ();
 sg13g2_fill_1 FILLER_4_2579 ();
 sg13g2_decap_8 FILLER_4_2593 ();
 sg13g2_decap_8 FILLER_4_2600 ();
 sg13g2_decap_8 FILLER_4_2607 ();
 sg13g2_decap_8 FILLER_4_2614 ();
 sg13g2_fill_2 FILLER_4_2621 ();
 sg13g2_fill_1 FILLER_4_2623 ();
 sg13g2_decap_8 FILLER_4_2650 ();
 sg13g2_decap_8 FILLER_4_2657 ();
 sg13g2_decap_4 FILLER_4_2664 ();
 sg13g2_fill_1 FILLER_4_2668 ();
 sg13g2_decap_8 FILLER_4_2682 ();
 sg13g2_decap_8 FILLER_4_2689 ();
 sg13g2_decap_4 FILLER_4_2696 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_4 FILLER_5_497 ();
 sg13g2_fill_2 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_506 ();
 sg13g2_decap_8 FILLER_5_513 ();
 sg13g2_decap_8 FILLER_5_520 ();
 sg13g2_decap_8 FILLER_5_527 ();
 sg13g2_decap_8 FILLER_5_534 ();
 sg13g2_decap_8 FILLER_5_541 ();
 sg13g2_decap_4 FILLER_5_548 ();
 sg13g2_decap_8 FILLER_5_573 ();
 sg13g2_decap_8 FILLER_5_580 ();
 sg13g2_decap_8 FILLER_5_587 ();
 sg13g2_decap_8 FILLER_5_594 ();
 sg13g2_decap_8 FILLER_5_601 ();
 sg13g2_decap_8 FILLER_5_608 ();
 sg13g2_decap_8 FILLER_5_615 ();
 sg13g2_fill_2 FILLER_5_622 ();
 sg13g2_decap_8 FILLER_5_666 ();
 sg13g2_decap_8 FILLER_5_673 ();
 sg13g2_decap_8 FILLER_5_680 ();
 sg13g2_decap_8 FILLER_5_687 ();
 sg13g2_decap_8 FILLER_5_694 ();
 sg13g2_decap_8 FILLER_5_701 ();
 sg13g2_decap_8 FILLER_5_708 ();
 sg13g2_decap_8 FILLER_5_715 ();
 sg13g2_decap_8 FILLER_5_722 ();
 sg13g2_decap_8 FILLER_5_729 ();
 sg13g2_decap_8 FILLER_5_736 ();
 sg13g2_decap_4 FILLER_5_743 ();
 sg13g2_fill_1 FILLER_5_747 ();
 sg13g2_decap_4 FILLER_5_773 ();
 sg13g2_fill_2 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_804 ();
 sg13g2_decap_8 FILLER_5_811 ();
 sg13g2_decap_8 FILLER_5_818 ();
 sg13g2_decap_8 FILLER_5_825 ();
 sg13g2_decap_8 FILLER_5_832 ();
 sg13g2_decap_8 FILLER_5_839 ();
 sg13g2_decap_8 FILLER_5_846 ();
 sg13g2_decap_8 FILLER_5_853 ();
 sg13g2_decap_8 FILLER_5_860 ();
 sg13g2_decap_8 FILLER_5_867 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_decap_8 FILLER_5_881 ();
 sg13g2_decap_8 FILLER_5_888 ();
 sg13g2_decap_8 FILLER_5_895 ();
 sg13g2_decap_8 FILLER_5_902 ();
 sg13g2_decap_8 FILLER_5_909 ();
 sg13g2_decap_8 FILLER_5_916 ();
 sg13g2_decap_8 FILLER_5_923 ();
 sg13g2_decap_8 FILLER_5_930 ();
 sg13g2_decap_8 FILLER_5_937 ();
 sg13g2_decap_8 FILLER_5_944 ();
 sg13g2_decap_8 FILLER_5_951 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_decap_8 FILLER_5_965 ();
 sg13g2_decap_8 FILLER_5_972 ();
 sg13g2_decap_8 FILLER_5_979 ();
 sg13g2_decap_8 FILLER_5_986 ();
 sg13g2_decap_8 FILLER_5_993 ();
 sg13g2_decap_8 FILLER_5_1000 ();
 sg13g2_decap_4 FILLER_5_1007 ();
 sg13g2_decap_8 FILLER_5_1032 ();
 sg13g2_decap_8 FILLER_5_1039 ();
 sg13g2_decap_4 FILLER_5_1046 ();
 sg13g2_decap_8 FILLER_5_1071 ();
 sg13g2_decap_8 FILLER_5_1078 ();
 sg13g2_decap_8 FILLER_5_1085 ();
 sg13g2_decap_8 FILLER_5_1092 ();
 sg13g2_decap_8 FILLER_5_1099 ();
 sg13g2_decap_8 FILLER_5_1106 ();
 sg13g2_decap_8 FILLER_5_1113 ();
 sg13g2_decap_8 FILLER_5_1120 ();
 sg13g2_decap_8 FILLER_5_1127 ();
 sg13g2_decap_8 FILLER_5_1134 ();
 sg13g2_decap_8 FILLER_5_1141 ();
 sg13g2_decap_8 FILLER_5_1148 ();
 sg13g2_decap_8 FILLER_5_1155 ();
 sg13g2_decap_8 FILLER_5_1162 ();
 sg13g2_decap_8 FILLER_5_1169 ();
 sg13g2_decap_8 FILLER_5_1176 ();
 sg13g2_decap_8 FILLER_5_1183 ();
 sg13g2_decap_8 FILLER_5_1190 ();
 sg13g2_decap_8 FILLER_5_1197 ();
 sg13g2_decap_8 FILLER_5_1204 ();
 sg13g2_fill_2 FILLER_5_1211 ();
 sg13g2_decap_8 FILLER_5_1234 ();
 sg13g2_decap_8 FILLER_5_1241 ();
 sg13g2_decap_4 FILLER_5_1248 ();
 sg13g2_fill_1 FILLER_5_1252 ();
 sg13g2_decap_8 FILLER_5_1278 ();
 sg13g2_decap_8 FILLER_5_1285 ();
 sg13g2_decap_8 FILLER_5_1292 ();
 sg13g2_fill_2 FILLER_5_1299 ();
 sg13g2_decap_8 FILLER_5_1326 ();
 sg13g2_decap_8 FILLER_5_1333 ();
 sg13g2_decap_8 FILLER_5_1340 ();
 sg13g2_decap_8 FILLER_5_1347 ();
 sg13g2_decap_8 FILLER_5_1354 ();
 sg13g2_decap_8 FILLER_5_1361 ();
 sg13g2_decap_8 FILLER_5_1368 ();
 sg13g2_decap_8 FILLER_5_1375 ();
 sg13g2_decap_8 FILLER_5_1382 ();
 sg13g2_decap_8 FILLER_5_1389 ();
 sg13g2_decap_8 FILLER_5_1396 ();
 sg13g2_decap_8 FILLER_5_1403 ();
 sg13g2_decap_8 FILLER_5_1410 ();
 sg13g2_decap_8 FILLER_5_1417 ();
 sg13g2_decap_4 FILLER_5_1424 ();
 sg13g2_fill_2 FILLER_5_1428 ();
 sg13g2_decap_8 FILLER_5_1433 ();
 sg13g2_decap_8 FILLER_5_1440 ();
 sg13g2_decap_8 FILLER_5_1447 ();
 sg13g2_decap_8 FILLER_5_1454 ();
 sg13g2_decap_8 FILLER_5_1461 ();
 sg13g2_decap_8 FILLER_5_1468 ();
 sg13g2_decap_8 FILLER_5_1475 ();
 sg13g2_fill_2 FILLER_5_1482 ();
 sg13g2_fill_1 FILLER_5_1484 ();
 sg13g2_decap_8 FILLER_5_1488 ();
 sg13g2_decap_8 FILLER_5_1495 ();
 sg13g2_decap_8 FILLER_5_1502 ();
 sg13g2_decap_8 FILLER_5_1509 ();
 sg13g2_decap_8 FILLER_5_1516 ();
 sg13g2_decap_8 FILLER_5_1523 ();
 sg13g2_decap_8 FILLER_5_1530 ();
 sg13g2_decap_8 FILLER_5_1537 ();
 sg13g2_decap_8 FILLER_5_1544 ();
 sg13g2_decap_8 FILLER_5_1551 ();
 sg13g2_decap_8 FILLER_5_1558 ();
 sg13g2_decap_8 FILLER_5_1565 ();
 sg13g2_decap_8 FILLER_5_1572 ();
 sg13g2_decap_8 FILLER_5_1579 ();
 sg13g2_decap_8 FILLER_5_1586 ();
 sg13g2_decap_8 FILLER_5_1593 ();
 sg13g2_decap_8 FILLER_5_1600 ();
 sg13g2_decap_8 FILLER_5_1607 ();
 sg13g2_decap_8 FILLER_5_1614 ();
 sg13g2_decap_8 FILLER_5_1621 ();
 sg13g2_decap_8 FILLER_5_1628 ();
 sg13g2_decap_8 FILLER_5_1635 ();
 sg13g2_decap_8 FILLER_5_1642 ();
 sg13g2_decap_8 FILLER_5_1649 ();
 sg13g2_decap_8 FILLER_5_1656 ();
 sg13g2_decap_8 FILLER_5_1663 ();
 sg13g2_decap_8 FILLER_5_1670 ();
 sg13g2_decap_8 FILLER_5_1677 ();
 sg13g2_decap_8 FILLER_5_1684 ();
 sg13g2_decap_8 FILLER_5_1691 ();
 sg13g2_decap_8 FILLER_5_1698 ();
 sg13g2_decap_8 FILLER_5_1705 ();
 sg13g2_decap_8 FILLER_5_1712 ();
 sg13g2_decap_8 FILLER_5_1719 ();
 sg13g2_decap_8 FILLER_5_1726 ();
 sg13g2_decap_8 FILLER_5_1733 ();
 sg13g2_decap_8 FILLER_5_1740 ();
 sg13g2_decap_8 FILLER_5_1747 ();
 sg13g2_decap_8 FILLER_5_1754 ();
 sg13g2_decap_8 FILLER_5_1761 ();
 sg13g2_decap_8 FILLER_5_1768 ();
 sg13g2_decap_8 FILLER_5_1775 ();
 sg13g2_decap_8 FILLER_5_1782 ();
 sg13g2_decap_8 FILLER_5_1789 ();
 sg13g2_decap_8 FILLER_5_1796 ();
 sg13g2_decap_8 FILLER_5_1803 ();
 sg13g2_decap_8 FILLER_5_1810 ();
 sg13g2_decap_8 FILLER_5_1817 ();
 sg13g2_decap_8 FILLER_5_1824 ();
 sg13g2_decap_8 FILLER_5_1831 ();
 sg13g2_decap_8 FILLER_5_1838 ();
 sg13g2_decap_8 FILLER_5_1845 ();
 sg13g2_decap_8 FILLER_5_1852 ();
 sg13g2_decap_8 FILLER_5_1859 ();
 sg13g2_decap_8 FILLER_5_1866 ();
 sg13g2_decap_8 FILLER_5_1873 ();
 sg13g2_decap_8 FILLER_5_1880 ();
 sg13g2_decap_8 FILLER_5_1887 ();
 sg13g2_decap_8 FILLER_5_1894 ();
 sg13g2_decap_8 FILLER_5_1901 ();
 sg13g2_decap_8 FILLER_5_1908 ();
 sg13g2_fill_1 FILLER_5_1915 ();
 sg13g2_decap_8 FILLER_5_1937 ();
 sg13g2_decap_8 FILLER_5_1944 ();
 sg13g2_decap_8 FILLER_5_1951 ();
 sg13g2_decap_8 FILLER_5_1958 ();
 sg13g2_decap_8 FILLER_5_1965 ();
 sg13g2_decap_8 FILLER_5_1972 ();
 sg13g2_decap_8 FILLER_5_1979 ();
 sg13g2_decap_8 FILLER_5_1986 ();
 sg13g2_decap_8 FILLER_5_1993 ();
 sg13g2_decap_8 FILLER_5_2000 ();
 sg13g2_decap_8 FILLER_5_2007 ();
 sg13g2_decap_8 FILLER_5_2014 ();
 sg13g2_decap_8 FILLER_5_2021 ();
 sg13g2_decap_8 FILLER_5_2028 ();
 sg13g2_decap_8 FILLER_5_2035 ();
 sg13g2_decap_8 FILLER_5_2042 ();
 sg13g2_decap_8 FILLER_5_2049 ();
 sg13g2_decap_8 FILLER_5_2056 ();
 sg13g2_decap_8 FILLER_5_2063 ();
 sg13g2_decap_8 FILLER_5_2070 ();
 sg13g2_decap_8 FILLER_5_2077 ();
 sg13g2_decap_8 FILLER_5_2084 ();
 sg13g2_decap_8 FILLER_5_2091 ();
 sg13g2_decap_8 FILLER_5_2119 ();
 sg13g2_decap_8 FILLER_5_2126 ();
 sg13g2_decap_8 FILLER_5_2133 ();
 sg13g2_decap_8 FILLER_5_2140 ();
 sg13g2_decap_8 FILLER_5_2147 ();
 sg13g2_decap_8 FILLER_5_2154 ();
 sg13g2_decap_8 FILLER_5_2161 ();
 sg13g2_decap_8 FILLER_5_2193 ();
 sg13g2_decap_8 FILLER_5_2200 ();
 sg13g2_decap_4 FILLER_5_2207 ();
 sg13g2_decap_8 FILLER_5_2236 ();
 sg13g2_decap_8 FILLER_5_2243 ();
 sg13g2_decap_8 FILLER_5_2250 ();
 sg13g2_decap_4 FILLER_5_2257 ();
 sg13g2_decap_8 FILLER_5_2276 ();
 sg13g2_decap_8 FILLER_5_2283 ();
 sg13g2_decap_8 FILLER_5_2290 ();
 sg13g2_decap_8 FILLER_5_2297 ();
 sg13g2_fill_2 FILLER_5_2304 ();
 sg13g2_fill_1 FILLER_5_2306 ();
 sg13g2_fill_1 FILLER_5_2322 ();
 sg13g2_decap_8 FILLER_5_2338 ();
 sg13g2_fill_2 FILLER_5_2345 ();
 sg13g2_fill_1 FILLER_5_2347 ();
 sg13g2_decap_8 FILLER_5_2373 ();
 sg13g2_fill_2 FILLER_5_2380 ();
 sg13g2_fill_1 FILLER_5_2382 ();
 sg13g2_decap_8 FILLER_5_2408 ();
 sg13g2_fill_2 FILLER_5_2415 ();
 sg13g2_fill_1 FILLER_5_2417 ();
 sg13g2_decap_8 FILLER_5_2443 ();
 sg13g2_decap_8 FILLER_5_2450 ();
 sg13g2_decap_8 FILLER_5_2457 ();
 sg13g2_fill_2 FILLER_5_2464 ();
 sg13g2_fill_1 FILLER_5_2466 ();
 sg13g2_decap_8 FILLER_5_2472 ();
 sg13g2_decap_8 FILLER_5_2479 ();
 sg13g2_decap_8 FILLER_5_2486 ();
 sg13g2_decap_8 FILLER_5_2493 ();
 sg13g2_decap_4 FILLER_5_2500 ();
 sg13g2_fill_2 FILLER_5_2504 ();
 sg13g2_decap_8 FILLER_5_2511 ();
 sg13g2_decap_8 FILLER_5_2518 ();
 sg13g2_decap_8 FILLER_5_2525 ();
 sg13g2_decap_8 FILLER_5_2532 ();
 sg13g2_decap_8 FILLER_5_2544 ();
 sg13g2_decap_8 FILLER_5_2551 ();
 sg13g2_decap_4 FILLER_5_2558 ();
 sg13g2_fill_2 FILLER_5_2562 ();
 sg13g2_decap_8 FILLER_5_2577 ();
 sg13g2_decap_4 FILLER_5_2584 ();
 sg13g2_decap_4 FILLER_5_2594 ();
 sg13g2_decap_8 FILLER_5_2611 ();
 sg13g2_decap_8 FILLER_5_2618 ();
 sg13g2_decap_8 FILLER_5_2625 ();
 sg13g2_fill_1 FILLER_5_2632 ();
 sg13g2_decap_4 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2649 ();
 sg13g2_decap_8 FILLER_5_2656 ();
 sg13g2_decap_8 FILLER_5_2663 ();
 sg13g2_fill_2 FILLER_5_2670 ();
 sg13g2_fill_1 FILLER_5_2672 ();
 sg13g2_fill_2 FILLER_5_2679 ();
 sg13g2_decap_8 FILLER_5_2687 ();
 sg13g2_decap_4 FILLER_5_2694 ();
 sg13g2_fill_2 FILLER_5_2698 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_521 ();
 sg13g2_decap_8 FILLER_6_528 ();
 sg13g2_decap_8 FILLER_6_535 ();
 sg13g2_decap_8 FILLER_6_542 ();
 sg13g2_decap_8 FILLER_6_549 ();
 sg13g2_decap_8 FILLER_6_556 ();
 sg13g2_decap_8 FILLER_6_563 ();
 sg13g2_decap_8 FILLER_6_570 ();
 sg13g2_decap_8 FILLER_6_577 ();
 sg13g2_decap_8 FILLER_6_584 ();
 sg13g2_decap_8 FILLER_6_591 ();
 sg13g2_decap_8 FILLER_6_598 ();
 sg13g2_decap_8 FILLER_6_605 ();
 sg13g2_decap_8 FILLER_6_612 ();
 sg13g2_decap_8 FILLER_6_619 ();
 sg13g2_decap_8 FILLER_6_626 ();
 sg13g2_decap_8 FILLER_6_633 ();
 sg13g2_decap_8 FILLER_6_640 ();
 sg13g2_decap_8 FILLER_6_647 ();
 sg13g2_decap_8 FILLER_6_654 ();
 sg13g2_decap_8 FILLER_6_661 ();
 sg13g2_decap_8 FILLER_6_668 ();
 sg13g2_decap_8 FILLER_6_675 ();
 sg13g2_fill_2 FILLER_6_682 ();
 sg13g2_decap_8 FILLER_6_687 ();
 sg13g2_decap_8 FILLER_6_694 ();
 sg13g2_decap_8 FILLER_6_701 ();
 sg13g2_decap_8 FILLER_6_708 ();
 sg13g2_fill_1 FILLER_6_715 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_4 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_848 ();
 sg13g2_decap_8 FILLER_6_855 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_869 ();
 sg13g2_decap_8 FILLER_6_876 ();
 sg13g2_decap_8 FILLER_6_883 ();
 sg13g2_decap_8 FILLER_6_890 ();
 sg13g2_decap_8 FILLER_6_897 ();
 sg13g2_decap_8 FILLER_6_904 ();
 sg13g2_decap_8 FILLER_6_911 ();
 sg13g2_decap_8 FILLER_6_918 ();
 sg13g2_decap_8 FILLER_6_925 ();
 sg13g2_decap_8 FILLER_6_932 ();
 sg13g2_decap_8 FILLER_6_939 ();
 sg13g2_decap_8 FILLER_6_946 ();
 sg13g2_decap_8 FILLER_6_953 ();
 sg13g2_decap_8 FILLER_6_960 ();
 sg13g2_decap_8 FILLER_6_967 ();
 sg13g2_decap_8 FILLER_6_974 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_fill_1 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1031 ();
 sg13g2_decap_8 FILLER_6_1038 ();
 sg13g2_fill_2 FILLER_6_1045 ();
 sg13g2_fill_1 FILLER_6_1047 ();
 sg13g2_decap_8 FILLER_6_1073 ();
 sg13g2_decap_8 FILLER_6_1080 ();
 sg13g2_decap_8 FILLER_6_1087 ();
 sg13g2_decap_4 FILLER_6_1094 ();
 sg13g2_decap_8 FILLER_6_1119 ();
 sg13g2_decap_8 FILLER_6_1126 ();
 sg13g2_decap_8 FILLER_6_1133 ();
 sg13g2_decap_8 FILLER_6_1140 ();
 sg13g2_decap_8 FILLER_6_1147 ();
 sg13g2_decap_8 FILLER_6_1154 ();
 sg13g2_decap_8 FILLER_6_1161 ();
 sg13g2_decap_8 FILLER_6_1168 ();
 sg13g2_decap_8 FILLER_6_1175 ();
 sg13g2_decap_8 FILLER_6_1182 ();
 sg13g2_decap_8 FILLER_6_1189 ();
 sg13g2_decap_8 FILLER_6_1196 ();
 sg13g2_decap_8 FILLER_6_1203 ();
 sg13g2_decap_8 FILLER_6_1235 ();
 sg13g2_decap_8 FILLER_6_1242 ();
 sg13g2_decap_8 FILLER_6_1249 ();
 sg13g2_decap_8 FILLER_6_1256 ();
 sg13g2_decap_8 FILLER_6_1263 ();
 sg13g2_decap_8 FILLER_6_1270 ();
 sg13g2_decap_8 FILLER_6_1277 ();
 sg13g2_decap_8 FILLER_6_1284 ();
 sg13g2_decap_8 FILLER_6_1291 ();
 sg13g2_decap_8 FILLER_6_1298 ();
 sg13g2_decap_8 FILLER_6_1305 ();
 sg13g2_decap_8 FILLER_6_1312 ();
 sg13g2_decap_8 FILLER_6_1319 ();
 sg13g2_decap_8 FILLER_6_1326 ();
 sg13g2_decap_8 FILLER_6_1333 ();
 sg13g2_decap_8 FILLER_6_1340 ();
 sg13g2_decap_8 FILLER_6_1347 ();
 sg13g2_decap_8 FILLER_6_1354 ();
 sg13g2_decap_8 FILLER_6_1361 ();
 sg13g2_decap_8 FILLER_6_1368 ();
 sg13g2_decap_8 FILLER_6_1375 ();
 sg13g2_decap_8 FILLER_6_1382 ();
 sg13g2_decap_8 FILLER_6_1389 ();
 sg13g2_decap_8 FILLER_6_1396 ();
 sg13g2_decap_8 FILLER_6_1403 ();
 sg13g2_decap_8 FILLER_6_1410 ();
 sg13g2_decap_8 FILLER_6_1417 ();
 sg13g2_decap_8 FILLER_6_1424 ();
 sg13g2_decap_8 FILLER_6_1431 ();
 sg13g2_decap_8 FILLER_6_1438 ();
 sg13g2_decap_8 FILLER_6_1445 ();
 sg13g2_decap_8 FILLER_6_1452 ();
 sg13g2_decap_8 FILLER_6_1459 ();
 sg13g2_decap_8 FILLER_6_1466 ();
 sg13g2_decap_8 FILLER_6_1473 ();
 sg13g2_decap_8 FILLER_6_1480 ();
 sg13g2_decap_4 FILLER_6_1487 ();
 sg13g2_fill_1 FILLER_6_1491 ();
 sg13g2_decap_8 FILLER_6_1495 ();
 sg13g2_decap_8 FILLER_6_1502 ();
 sg13g2_decap_8 FILLER_6_1509 ();
 sg13g2_decap_8 FILLER_6_1516 ();
 sg13g2_decap_8 FILLER_6_1523 ();
 sg13g2_decap_8 FILLER_6_1530 ();
 sg13g2_decap_8 FILLER_6_1537 ();
 sg13g2_decap_8 FILLER_6_1544 ();
 sg13g2_decap_8 FILLER_6_1551 ();
 sg13g2_decap_8 FILLER_6_1558 ();
 sg13g2_decap_8 FILLER_6_1565 ();
 sg13g2_fill_1 FILLER_6_1572 ();
 sg13g2_decap_8 FILLER_6_1576 ();
 sg13g2_decap_8 FILLER_6_1583 ();
 sg13g2_decap_8 FILLER_6_1590 ();
 sg13g2_decap_8 FILLER_6_1597 ();
 sg13g2_decap_8 FILLER_6_1604 ();
 sg13g2_decap_8 FILLER_6_1611 ();
 sg13g2_decap_8 FILLER_6_1618 ();
 sg13g2_decap_8 FILLER_6_1625 ();
 sg13g2_decap_8 FILLER_6_1632 ();
 sg13g2_decap_8 FILLER_6_1639 ();
 sg13g2_decap_8 FILLER_6_1646 ();
 sg13g2_decap_8 FILLER_6_1653 ();
 sg13g2_decap_8 FILLER_6_1660 ();
 sg13g2_decap_8 FILLER_6_1667 ();
 sg13g2_decap_8 FILLER_6_1674 ();
 sg13g2_decap_8 FILLER_6_1681 ();
 sg13g2_decap_8 FILLER_6_1688 ();
 sg13g2_decap_8 FILLER_6_1695 ();
 sg13g2_decap_8 FILLER_6_1702 ();
 sg13g2_decap_8 FILLER_6_1709 ();
 sg13g2_decap_8 FILLER_6_1716 ();
 sg13g2_decap_8 FILLER_6_1723 ();
 sg13g2_decap_8 FILLER_6_1730 ();
 sg13g2_decap_8 FILLER_6_1737 ();
 sg13g2_decap_8 FILLER_6_1744 ();
 sg13g2_decap_8 FILLER_6_1751 ();
 sg13g2_decap_8 FILLER_6_1758 ();
 sg13g2_decap_8 FILLER_6_1765 ();
 sg13g2_decap_8 FILLER_6_1772 ();
 sg13g2_decap_8 FILLER_6_1779 ();
 sg13g2_decap_8 FILLER_6_1786 ();
 sg13g2_decap_8 FILLER_6_1793 ();
 sg13g2_decap_8 FILLER_6_1800 ();
 sg13g2_decap_8 FILLER_6_1807 ();
 sg13g2_decap_8 FILLER_6_1814 ();
 sg13g2_decap_8 FILLER_6_1821 ();
 sg13g2_decap_8 FILLER_6_1828 ();
 sg13g2_decap_8 FILLER_6_1835 ();
 sg13g2_decap_8 FILLER_6_1842 ();
 sg13g2_decap_8 FILLER_6_1849 ();
 sg13g2_decap_8 FILLER_6_1856 ();
 sg13g2_decap_8 FILLER_6_1863 ();
 sg13g2_decap_8 FILLER_6_1870 ();
 sg13g2_decap_8 FILLER_6_1877 ();
 sg13g2_decap_8 FILLER_6_1884 ();
 sg13g2_decap_8 FILLER_6_1891 ();
 sg13g2_decap_8 FILLER_6_1898 ();
 sg13g2_decap_8 FILLER_6_1905 ();
 sg13g2_fill_2 FILLER_6_1912 ();
 sg13g2_decap_8 FILLER_6_1939 ();
 sg13g2_decap_8 FILLER_6_1946 ();
 sg13g2_decap_8 FILLER_6_1953 ();
 sg13g2_fill_1 FILLER_6_1960 ();
 sg13g2_decap_8 FILLER_6_1982 ();
 sg13g2_decap_8 FILLER_6_1989 ();
 sg13g2_decap_8 FILLER_6_1996 ();
 sg13g2_decap_8 FILLER_6_2003 ();
 sg13g2_decap_8 FILLER_6_2031 ();
 sg13g2_decap_8 FILLER_6_2038 ();
 sg13g2_decap_8 FILLER_6_2045 ();
 sg13g2_decap_8 FILLER_6_2052 ();
 sg13g2_decap_8 FILLER_6_2059 ();
 sg13g2_decap_8 FILLER_6_2066 ();
 sg13g2_decap_8 FILLER_6_2073 ();
 sg13g2_decap_8 FILLER_6_2080 ();
 sg13g2_decap_8 FILLER_6_2087 ();
 sg13g2_fill_1 FILLER_6_2094 ();
 sg13g2_decap_8 FILLER_6_2120 ();
 sg13g2_decap_8 FILLER_6_2127 ();
 sg13g2_decap_8 FILLER_6_2155 ();
 sg13g2_decap_8 FILLER_6_2162 ();
 sg13g2_decap_8 FILLER_6_2169 ();
 sg13g2_decap_8 FILLER_6_2176 ();
 sg13g2_decap_8 FILLER_6_2183 ();
 sg13g2_decap_8 FILLER_6_2190 ();
 sg13g2_decap_8 FILLER_6_2197 ();
 sg13g2_decap_8 FILLER_6_2204 ();
 sg13g2_decap_8 FILLER_6_2211 ();
 sg13g2_decap_8 FILLER_6_2218 ();
 sg13g2_decap_8 FILLER_6_2225 ();
 sg13g2_decap_8 FILLER_6_2232 ();
 sg13g2_decap_8 FILLER_6_2239 ();
 sg13g2_decap_8 FILLER_6_2246 ();
 sg13g2_decap_8 FILLER_6_2253 ();
 sg13g2_decap_4 FILLER_6_2260 ();
 sg13g2_fill_2 FILLER_6_2264 ();
 sg13g2_decap_8 FILLER_6_2281 ();
 sg13g2_decap_8 FILLER_6_2288 ();
 sg13g2_fill_2 FILLER_6_2295 ();
 sg13g2_fill_1 FILLER_6_2297 ();
 sg13g2_decap_8 FILLER_6_2313 ();
 sg13g2_decap_8 FILLER_6_2320 ();
 sg13g2_decap_8 FILLER_6_2327 ();
 sg13g2_decap_8 FILLER_6_2334 ();
 sg13g2_decap_8 FILLER_6_2341 ();
 sg13g2_decap_8 FILLER_6_2348 ();
 sg13g2_decap_8 FILLER_6_2355 ();
 sg13g2_decap_8 FILLER_6_2362 ();
 sg13g2_decap_8 FILLER_6_2369 ();
 sg13g2_decap_8 FILLER_6_2376 ();
 sg13g2_decap_8 FILLER_6_2383 ();
 sg13g2_decap_4 FILLER_6_2390 ();
 sg13g2_decap_8 FILLER_6_2399 ();
 sg13g2_decap_8 FILLER_6_2406 ();
 sg13g2_decap_8 FILLER_6_2413 ();
 sg13g2_decap_8 FILLER_6_2420 ();
 sg13g2_decap_8 FILLER_6_2427 ();
 sg13g2_decap_8 FILLER_6_2434 ();
 sg13g2_decap_8 FILLER_6_2441 ();
 sg13g2_decap_8 FILLER_6_2448 ();
 sg13g2_fill_1 FILLER_6_2455 ();
 sg13g2_decap_8 FILLER_6_2481 ();
 sg13g2_decap_8 FILLER_6_2488 ();
 sg13g2_decap_8 FILLER_6_2520 ();
 sg13g2_decap_8 FILLER_6_2527 ();
 sg13g2_decap_8 FILLER_6_2534 ();
 sg13g2_decap_8 FILLER_6_2541 ();
 sg13g2_decap_8 FILLER_6_2548 ();
 sg13g2_decap_8 FILLER_6_2555 ();
 sg13g2_decap_8 FILLER_6_2562 ();
 sg13g2_decap_4 FILLER_6_2569 ();
 sg13g2_fill_1 FILLER_6_2573 ();
 sg13g2_decap_8 FILLER_6_2580 ();
 sg13g2_decap_8 FILLER_6_2587 ();
 sg13g2_fill_2 FILLER_6_2594 ();
 sg13g2_fill_1 FILLER_6_2596 ();
 sg13g2_decap_4 FILLER_6_2600 ();
 sg13g2_fill_1 FILLER_6_2604 ();
 sg13g2_decap_8 FILLER_6_2611 ();
 sg13g2_decap_8 FILLER_6_2618 ();
 sg13g2_decap_8 FILLER_6_2625 ();
 sg13g2_decap_8 FILLER_6_2632 ();
 sg13g2_decap_8 FILLER_6_2639 ();
 sg13g2_decap_8 FILLER_6_2646 ();
 sg13g2_decap_8 FILLER_6_2653 ();
 sg13g2_decap_8 FILLER_6_2660 ();
 sg13g2_decap_4 FILLER_6_2667 ();
 sg13g2_fill_1 FILLER_6_2671 ();
 sg13g2_decap_4 FILLER_6_2678 ();
 sg13g2_fill_2 FILLER_6_2682 ();
 sg13g2_decap_8 FILLER_6_2687 ();
 sg13g2_decap_4 FILLER_6_2694 ();
 sg13g2_fill_2 FILLER_6_2698 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_fill_2 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_548 ();
 sg13g2_decap_8 FILLER_7_555 ();
 sg13g2_decap_8 FILLER_7_562 ();
 sg13g2_decap_8 FILLER_7_569 ();
 sg13g2_decap_4 FILLER_7_576 ();
 sg13g2_fill_1 FILLER_7_580 ();
 sg13g2_fill_2 FILLER_7_602 ();
 sg13g2_fill_1 FILLER_7_604 ();
 sg13g2_decap_8 FILLER_7_626 ();
 sg13g2_decap_8 FILLER_7_633 ();
 sg13g2_decap_8 FILLER_7_640 ();
 sg13g2_decap_8 FILLER_7_647 ();
 sg13g2_decap_8 FILLER_7_654 ();
 sg13g2_decap_8 FILLER_7_661 ();
 sg13g2_decap_8 FILLER_7_668 ();
 sg13g2_decap_8 FILLER_7_675 ();
 sg13g2_decap_8 FILLER_7_682 ();
 sg13g2_decap_8 FILLER_7_689 ();
 sg13g2_decap_8 FILLER_7_696 ();
 sg13g2_decap_4 FILLER_7_703 ();
 sg13g2_fill_1 FILLER_7_707 ();
 sg13g2_decap_4 FILLER_7_711 ();
 sg13g2_decap_8 FILLER_7_718 ();
 sg13g2_decap_8 FILLER_7_725 ();
 sg13g2_fill_1 FILLER_7_732 ();
 sg13g2_decap_8 FILLER_7_738 ();
 sg13g2_decap_8 FILLER_7_745 ();
 sg13g2_decap_8 FILLER_7_752 ();
 sg13g2_decap_8 FILLER_7_759 ();
 sg13g2_decap_8 FILLER_7_766 ();
 sg13g2_decap_8 FILLER_7_773 ();
 sg13g2_decap_8 FILLER_7_780 ();
 sg13g2_decap_8 FILLER_7_787 ();
 sg13g2_decap_8 FILLER_7_794 ();
 sg13g2_decap_8 FILLER_7_801 ();
 sg13g2_decap_8 FILLER_7_808 ();
 sg13g2_decap_8 FILLER_7_815 ();
 sg13g2_decap_8 FILLER_7_822 ();
 sg13g2_decap_8 FILLER_7_829 ();
 sg13g2_decap_8 FILLER_7_836 ();
 sg13g2_decap_8 FILLER_7_843 ();
 sg13g2_decap_8 FILLER_7_850 ();
 sg13g2_fill_2 FILLER_7_857 ();
 sg13g2_decap_8 FILLER_7_884 ();
 sg13g2_decap_4 FILLER_7_891 ();
 sg13g2_decap_8 FILLER_7_920 ();
 sg13g2_decap_8 FILLER_7_927 ();
 sg13g2_decap_8 FILLER_7_934 ();
 sg13g2_fill_1 FILLER_7_941 ();
 sg13g2_decap_8 FILLER_7_967 ();
 sg13g2_decap_8 FILLER_7_974 ();
 sg13g2_decap_8 FILLER_7_981 ();
 sg13g2_decap_8 FILLER_7_988 ();
 sg13g2_decap_8 FILLER_7_995 ();
 sg13g2_decap_8 FILLER_7_1002 ();
 sg13g2_decap_8 FILLER_7_1009 ();
 sg13g2_decap_8 FILLER_7_1016 ();
 sg13g2_decap_8 FILLER_7_1023 ();
 sg13g2_decap_8 FILLER_7_1030 ();
 sg13g2_decap_8 FILLER_7_1037 ();
 sg13g2_decap_8 FILLER_7_1044 ();
 sg13g2_decap_8 FILLER_7_1051 ();
 sg13g2_decap_8 FILLER_7_1058 ();
 sg13g2_decap_8 FILLER_7_1065 ();
 sg13g2_decap_8 FILLER_7_1072 ();
 sg13g2_decap_8 FILLER_7_1079 ();
 sg13g2_decap_4 FILLER_7_1086 ();
 sg13g2_decap_8 FILLER_7_1115 ();
 sg13g2_decap_8 FILLER_7_1122 ();
 sg13g2_decap_8 FILLER_7_1129 ();
 sg13g2_decap_8 FILLER_7_1136 ();
 sg13g2_decap_8 FILLER_7_1143 ();
 sg13g2_decap_8 FILLER_7_1150 ();
 sg13g2_decap_8 FILLER_7_1157 ();
 sg13g2_decap_8 FILLER_7_1164 ();
 sg13g2_decap_8 FILLER_7_1171 ();
 sg13g2_decap_8 FILLER_7_1178 ();
 sg13g2_decap_8 FILLER_7_1185 ();
 sg13g2_decap_8 FILLER_7_1192 ();
 sg13g2_decap_8 FILLER_7_1199 ();
 sg13g2_decap_8 FILLER_7_1206 ();
 sg13g2_decap_8 FILLER_7_1213 ();
 sg13g2_decap_8 FILLER_7_1220 ();
 sg13g2_decap_8 FILLER_7_1227 ();
 sg13g2_decap_8 FILLER_7_1234 ();
 sg13g2_decap_8 FILLER_7_1241 ();
 sg13g2_decap_8 FILLER_7_1248 ();
 sg13g2_decap_8 FILLER_7_1255 ();
 sg13g2_decap_8 FILLER_7_1262 ();
 sg13g2_decap_8 FILLER_7_1269 ();
 sg13g2_decap_8 FILLER_7_1276 ();
 sg13g2_decap_8 FILLER_7_1283 ();
 sg13g2_decap_8 FILLER_7_1290 ();
 sg13g2_decap_8 FILLER_7_1297 ();
 sg13g2_decap_8 FILLER_7_1304 ();
 sg13g2_decap_8 FILLER_7_1311 ();
 sg13g2_decap_8 FILLER_7_1318 ();
 sg13g2_decap_8 FILLER_7_1325 ();
 sg13g2_decap_8 FILLER_7_1332 ();
 sg13g2_decap_8 FILLER_7_1339 ();
 sg13g2_decap_8 FILLER_7_1346 ();
 sg13g2_decap_8 FILLER_7_1353 ();
 sg13g2_decap_8 FILLER_7_1360 ();
 sg13g2_decap_8 FILLER_7_1367 ();
 sg13g2_decap_8 FILLER_7_1374 ();
 sg13g2_decap_8 FILLER_7_1381 ();
 sg13g2_decap_8 FILLER_7_1388 ();
 sg13g2_decap_8 FILLER_7_1395 ();
 sg13g2_decap_8 FILLER_7_1402 ();
 sg13g2_decap_8 FILLER_7_1409 ();
 sg13g2_decap_8 FILLER_7_1416 ();
 sg13g2_decap_8 FILLER_7_1423 ();
 sg13g2_decap_8 FILLER_7_1430 ();
 sg13g2_decap_8 FILLER_7_1437 ();
 sg13g2_decap_8 FILLER_7_1444 ();
 sg13g2_decap_8 FILLER_7_1451 ();
 sg13g2_decap_8 FILLER_7_1458 ();
 sg13g2_decap_8 FILLER_7_1465 ();
 sg13g2_decap_8 FILLER_7_1472 ();
 sg13g2_decap_8 FILLER_7_1479 ();
 sg13g2_decap_8 FILLER_7_1486 ();
 sg13g2_decap_8 FILLER_7_1493 ();
 sg13g2_decap_8 FILLER_7_1500 ();
 sg13g2_fill_2 FILLER_7_1507 ();
 sg13g2_fill_1 FILLER_7_1509 ();
 sg13g2_decap_8 FILLER_7_1513 ();
 sg13g2_decap_8 FILLER_7_1520 ();
 sg13g2_decap_8 FILLER_7_1527 ();
 sg13g2_decap_8 FILLER_7_1534 ();
 sg13g2_decap_8 FILLER_7_1541 ();
 sg13g2_decap_8 FILLER_7_1548 ();
 sg13g2_decap_8 FILLER_7_1555 ();
 sg13g2_decap_8 FILLER_7_1562 ();
 sg13g2_decap_8 FILLER_7_1569 ();
 sg13g2_decap_8 FILLER_7_1576 ();
 sg13g2_decap_8 FILLER_7_1583 ();
 sg13g2_decap_8 FILLER_7_1590 ();
 sg13g2_decap_8 FILLER_7_1597 ();
 sg13g2_decap_8 FILLER_7_1604 ();
 sg13g2_decap_8 FILLER_7_1611 ();
 sg13g2_decap_8 FILLER_7_1618 ();
 sg13g2_decap_8 FILLER_7_1625 ();
 sg13g2_decap_8 FILLER_7_1632 ();
 sg13g2_decap_8 FILLER_7_1639 ();
 sg13g2_decap_8 FILLER_7_1646 ();
 sg13g2_decap_8 FILLER_7_1653 ();
 sg13g2_decap_8 FILLER_7_1660 ();
 sg13g2_decap_8 FILLER_7_1667 ();
 sg13g2_decap_8 FILLER_7_1674 ();
 sg13g2_decap_8 FILLER_7_1681 ();
 sg13g2_decap_8 FILLER_7_1688 ();
 sg13g2_decap_8 FILLER_7_1695 ();
 sg13g2_decap_8 FILLER_7_1702 ();
 sg13g2_decap_8 FILLER_7_1709 ();
 sg13g2_decap_8 FILLER_7_1716 ();
 sg13g2_decap_8 FILLER_7_1723 ();
 sg13g2_decap_8 FILLER_7_1730 ();
 sg13g2_decap_8 FILLER_7_1737 ();
 sg13g2_decap_8 FILLER_7_1744 ();
 sg13g2_decap_8 FILLER_7_1751 ();
 sg13g2_decap_8 FILLER_7_1758 ();
 sg13g2_decap_8 FILLER_7_1765 ();
 sg13g2_decap_8 FILLER_7_1772 ();
 sg13g2_decap_8 FILLER_7_1779 ();
 sg13g2_decap_8 FILLER_7_1786 ();
 sg13g2_decap_8 FILLER_7_1793 ();
 sg13g2_decap_8 FILLER_7_1800 ();
 sg13g2_decap_8 FILLER_7_1807 ();
 sg13g2_decap_8 FILLER_7_1814 ();
 sg13g2_decap_8 FILLER_7_1821 ();
 sg13g2_decap_8 FILLER_7_1828 ();
 sg13g2_decap_8 FILLER_7_1835 ();
 sg13g2_decap_8 FILLER_7_1842 ();
 sg13g2_decap_8 FILLER_7_1849 ();
 sg13g2_decap_8 FILLER_7_1856 ();
 sg13g2_decap_8 FILLER_7_1863 ();
 sg13g2_decap_8 FILLER_7_1870 ();
 sg13g2_decap_8 FILLER_7_1877 ();
 sg13g2_decap_8 FILLER_7_1884 ();
 sg13g2_decap_8 FILLER_7_1891 ();
 sg13g2_decap_8 FILLER_7_1898 ();
 sg13g2_decap_8 FILLER_7_1905 ();
 sg13g2_decap_8 FILLER_7_1912 ();
 sg13g2_decap_8 FILLER_7_1919 ();
 sg13g2_decap_8 FILLER_7_1926 ();
 sg13g2_decap_8 FILLER_7_1933 ();
 sg13g2_decap_8 FILLER_7_1940 ();
 sg13g2_decap_8 FILLER_7_1947 ();
 sg13g2_decap_4 FILLER_7_1954 ();
 sg13g2_fill_1 FILLER_7_1958 ();
 sg13g2_decap_8 FILLER_7_1984 ();
 sg13g2_decap_8 FILLER_7_1991 ();
 sg13g2_decap_8 FILLER_7_1998 ();
 sg13g2_fill_1 FILLER_7_2005 ();
 sg13g2_decap_8 FILLER_7_2031 ();
 sg13g2_decap_8 FILLER_7_2038 ();
 sg13g2_decap_8 FILLER_7_2045 ();
 sg13g2_decap_8 FILLER_7_2052 ();
 sg13g2_decap_8 FILLER_7_2059 ();
 sg13g2_decap_8 FILLER_7_2066 ();
 sg13g2_decap_8 FILLER_7_2073 ();
 sg13g2_decap_8 FILLER_7_2080 ();
 sg13g2_decap_8 FILLER_7_2087 ();
 sg13g2_decap_8 FILLER_7_2094 ();
 sg13g2_decap_8 FILLER_7_2101 ();
 sg13g2_decap_8 FILLER_7_2108 ();
 sg13g2_decap_8 FILLER_7_2115 ();
 sg13g2_decap_8 FILLER_7_2122 ();
 sg13g2_fill_2 FILLER_7_2129 ();
 sg13g2_decap_8 FILLER_7_2156 ();
 sg13g2_decap_8 FILLER_7_2163 ();
 sg13g2_decap_8 FILLER_7_2170 ();
 sg13g2_decap_8 FILLER_7_2177 ();
 sg13g2_decap_8 FILLER_7_2184 ();
 sg13g2_decap_8 FILLER_7_2191 ();
 sg13g2_decap_8 FILLER_7_2198 ();
 sg13g2_decap_8 FILLER_7_2205 ();
 sg13g2_decap_8 FILLER_7_2212 ();
 sg13g2_decap_8 FILLER_7_2219 ();
 sg13g2_decap_8 FILLER_7_2226 ();
 sg13g2_decap_8 FILLER_7_2233 ();
 sg13g2_decap_8 FILLER_7_2240 ();
 sg13g2_decap_8 FILLER_7_2247 ();
 sg13g2_decap_8 FILLER_7_2254 ();
 sg13g2_fill_2 FILLER_7_2261 ();
 sg13g2_decap_8 FILLER_7_2278 ();
 sg13g2_decap_8 FILLER_7_2285 ();
 sg13g2_decap_8 FILLER_7_2292 ();
 sg13g2_decap_8 FILLER_7_2299 ();
 sg13g2_decap_8 FILLER_7_2306 ();
 sg13g2_decap_8 FILLER_7_2313 ();
 sg13g2_decap_8 FILLER_7_2320 ();
 sg13g2_decap_8 FILLER_7_2327 ();
 sg13g2_decap_8 FILLER_7_2334 ();
 sg13g2_decap_4 FILLER_7_2341 ();
 sg13g2_decap_8 FILLER_7_2350 ();
 sg13g2_decap_8 FILLER_7_2357 ();
 sg13g2_decap_8 FILLER_7_2364 ();
 sg13g2_decap_8 FILLER_7_2371 ();
 sg13g2_decap_8 FILLER_7_2378 ();
 sg13g2_decap_8 FILLER_7_2385 ();
 sg13g2_decap_8 FILLER_7_2397 ();
 sg13g2_decap_8 FILLER_7_2404 ();
 sg13g2_decap_8 FILLER_7_2411 ();
 sg13g2_decap_8 FILLER_7_2418 ();
 sg13g2_decap_8 FILLER_7_2425 ();
 sg13g2_fill_1 FILLER_7_2432 ();
 sg13g2_decap_8 FILLER_7_2438 ();
 sg13g2_decap_8 FILLER_7_2445 ();
 sg13g2_decap_8 FILLER_7_2452 ();
 sg13g2_decap_8 FILLER_7_2459 ();
 sg13g2_decap_8 FILLER_7_2466 ();
 sg13g2_decap_8 FILLER_7_2473 ();
 sg13g2_decap_8 FILLER_7_2480 ();
 sg13g2_decap_8 FILLER_7_2487 ();
 sg13g2_decap_8 FILLER_7_2494 ();
 sg13g2_decap_8 FILLER_7_2501 ();
 sg13g2_decap_8 FILLER_7_2508 ();
 sg13g2_decap_8 FILLER_7_2515 ();
 sg13g2_decap_8 FILLER_7_2522 ();
 sg13g2_decap_8 FILLER_7_2529 ();
 sg13g2_decap_8 FILLER_7_2536 ();
 sg13g2_decap_4 FILLER_7_2543 ();
 sg13g2_fill_1 FILLER_7_2547 ();
 sg13g2_fill_2 FILLER_7_2554 ();
 sg13g2_decap_8 FILLER_7_2562 ();
 sg13g2_decap_8 FILLER_7_2569 ();
 sg13g2_decap_8 FILLER_7_2576 ();
 sg13g2_fill_2 FILLER_7_2583 ();
 sg13g2_decap_8 FILLER_7_2588 ();
 sg13g2_decap_8 FILLER_7_2595 ();
 sg13g2_decap_8 FILLER_7_2602 ();
 sg13g2_decap_4 FILLER_7_2609 ();
 sg13g2_fill_1 FILLER_7_2613 ();
 sg13g2_decap_8 FILLER_7_2617 ();
 sg13g2_decap_8 FILLER_7_2624 ();
 sg13g2_decap_8 FILLER_7_2631 ();
 sg13g2_decap_8 FILLER_7_2638 ();
 sg13g2_decap_8 FILLER_7_2645 ();
 sg13g2_decap_8 FILLER_7_2652 ();
 sg13g2_decap_8 FILLER_7_2659 ();
 sg13g2_fill_1 FILLER_7_2666 ();
 sg13g2_fill_2 FILLER_7_2680 ();
 sg13g2_fill_1 FILLER_7_2682 ();
 sg13g2_decap_8 FILLER_7_2690 ();
 sg13g2_fill_2 FILLER_7_2697 ();
 sg13g2_fill_1 FILLER_7_2699 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_4 FILLER_8_630 ();
 sg13g2_fill_2 FILLER_8_634 ();
 sg13g2_decap_8 FILLER_8_657 ();
 sg13g2_decap_8 FILLER_8_664 ();
 sg13g2_decap_4 FILLER_8_671 ();
 sg13g2_fill_2 FILLER_8_675 ();
 sg13g2_decap_8 FILLER_8_698 ();
 sg13g2_fill_2 FILLER_8_705 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_4 FILLER_8_756 ();
 sg13g2_fill_2 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_787 ();
 sg13g2_fill_2 FILLER_8_794 ();
 sg13g2_decap_8 FILLER_8_821 ();
 sg13g2_decap_8 FILLER_8_828 ();
 sg13g2_decap_8 FILLER_8_835 ();
 sg13g2_decap_8 FILLER_8_842 ();
 sg13g2_decap_8 FILLER_8_849 ();
 sg13g2_decap_8 FILLER_8_856 ();
 sg13g2_decap_8 FILLER_8_863 ();
 sg13g2_decap_8 FILLER_8_870 ();
 sg13g2_decap_8 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_8_884 ();
 sg13g2_decap_8 FILLER_8_891 ();
 sg13g2_decap_8 FILLER_8_898 ();
 sg13g2_decap_8 FILLER_8_905 ();
 sg13g2_decap_8 FILLER_8_912 ();
 sg13g2_decap_8 FILLER_8_919 ();
 sg13g2_decap_8 FILLER_8_926 ();
 sg13g2_decap_8 FILLER_8_958 ();
 sg13g2_decap_8 FILLER_8_965 ();
 sg13g2_decap_8 FILLER_8_972 ();
 sg13g2_decap_8 FILLER_8_979 ();
 sg13g2_decap_8 FILLER_8_986 ();
 sg13g2_decap_8 FILLER_8_993 ();
 sg13g2_decap_8 FILLER_8_1000 ();
 sg13g2_decap_8 FILLER_8_1007 ();
 sg13g2_decap_8 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1021 ();
 sg13g2_decap_8 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_8_1035 ();
 sg13g2_decap_8 FILLER_8_1042 ();
 sg13g2_decap_8 FILLER_8_1049 ();
 sg13g2_decap_8 FILLER_8_1056 ();
 sg13g2_decap_8 FILLER_8_1063 ();
 sg13g2_decap_8 FILLER_8_1070 ();
 sg13g2_decap_8 FILLER_8_1077 ();
 sg13g2_decap_8 FILLER_8_1084 ();
 sg13g2_decap_8 FILLER_8_1091 ();
 sg13g2_decap_8 FILLER_8_1098 ();
 sg13g2_decap_8 FILLER_8_1105 ();
 sg13g2_decap_8 FILLER_8_1112 ();
 sg13g2_decap_8 FILLER_8_1119 ();
 sg13g2_decap_4 FILLER_8_1126 ();
 sg13g2_fill_2 FILLER_8_1130 ();
 sg13g2_decap_8 FILLER_8_1153 ();
 sg13g2_decap_8 FILLER_8_1160 ();
 sg13g2_fill_2 FILLER_8_1167 ();
 sg13g2_fill_1 FILLER_8_1169 ();
 sg13g2_decap_8 FILLER_8_1195 ();
 sg13g2_decap_8 FILLER_8_1202 ();
 sg13g2_decap_8 FILLER_8_1209 ();
 sg13g2_decap_8 FILLER_8_1216 ();
 sg13g2_decap_8 FILLER_8_1223 ();
 sg13g2_decap_8 FILLER_8_1230 ();
 sg13g2_decap_8 FILLER_8_1237 ();
 sg13g2_decap_8 FILLER_8_1244 ();
 sg13g2_decap_4 FILLER_8_1251 ();
 sg13g2_decap_8 FILLER_8_1276 ();
 sg13g2_decap_8 FILLER_8_1283 ();
 sg13g2_decap_8 FILLER_8_1290 ();
 sg13g2_decap_4 FILLER_8_1297 ();
 sg13g2_decap_8 FILLER_8_1322 ();
 sg13g2_decap_8 FILLER_8_1329 ();
 sg13g2_decap_8 FILLER_8_1336 ();
 sg13g2_decap_8 FILLER_8_1343 ();
 sg13g2_decap_8 FILLER_8_1350 ();
 sg13g2_decap_8 FILLER_8_1357 ();
 sg13g2_decap_8 FILLER_8_1364 ();
 sg13g2_decap_8 FILLER_8_1371 ();
 sg13g2_decap_8 FILLER_8_1378 ();
 sg13g2_decap_8 FILLER_8_1385 ();
 sg13g2_decap_8 FILLER_8_1392 ();
 sg13g2_decap_8 FILLER_8_1399 ();
 sg13g2_decap_8 FILLER_8_1406 ();
 sg13g2_decap_8 FILLER_8_1413 ();
 sg13g2_decap_8 FILLER_8_1420 ();
 sg13g2_decap_8 FILLER_8_1427 ();
 sg13g2_decap_8 FILLER_8_1434 ();
 sg13g2_decap_8 FILLER_8_1441 ();
 sg13g2_decap_8 FILLER_8_1448 ();
 sg13g2_decap_8 FILLER_8_1455 ();
 sg13g2_decap_8 FILLER_8_1462 ();
 sg13g2_decap_8 FILLER_8_1469 ();
 sg13g2_decap_4 FILLER_8_1476 ();
 sg13g2_fill_2 FILLER_8_1480 ();
 sg13g2_decap_8 FILLER_8_1485 ();
 sg13g2_decap_8 FILLER_8_1492 ();
 sg13g2_decap_8 FILLER_8_1499 ();
 sg13g2_decap_8 FILLER_8_1506 ();
 sg13g2_decap_8 FILLER_8_1513 ();
 sg13g2_decap_8 FILLER_8_1520 ();
 sg13g2_decap_8 FILLER_8_1527 ();
 sg13g2_decap_8 FILLER_8_1534 ();
 sg13g2_decap_8 FILLER_8_1541 ();
 sg13g2_decap_8 FILLER_8_1548 ();
 sg13g2_fill_2 FILLER_8_1555 ();
 sg13g2_fill_1 FILLER_8_1557 ();
 sg13g2_decap_8 FILLER_8_1561 ();
 sg13g2_decap_8 FILLER_8_1568 ();
 sg13g2_decap_8 FILLER_8_1575 ();
 sg13g2_decap_8 FILLER_8_1582 ();
 sg13g2_decap_8 FILLER_8_1589 ();
 sg13g2_decap_8 FILLER_8_1596 ();
 sg13g2_decap_8 FILLER_8_1603 ();
 sg13g2_decap_8 FILLER_8_1610 ();
 sg13g2_decap_8 FILLER_8_1617 ();
 sg13g2_decap_8 FILLER_8_1624 ();
 sg13g2_decap_8 FILLER_8_1631 ();
 sg13g2_decap_8 FILLER_8_1638 ();
 sg13g2_decap_8 FILLER_8_1645 ();
 sg13g2_decap_8 FILLER_8_1652 ();
 sg13g2_decap_8 FILLER_8_1659 ();
 sg13g2_decap_8 FILLER_8_1666 ();
 sg13g2_decap_8 FILLER_8_1673 ();
 sg13g2_decap_8 FILLER_8_1680 ();
 sg13g2_decap_8 FILLER_8_1687 ();
 sg13g2_decap_8 FILLER_8_1694 ();
 sg13g2_decap_8 FILLER_8_1701 ();
 sg13g2_decap_8 FILLER_8_1708 ();
 sg13g2_decap_8 FILLER_8_1715 ();
 sg13g2_decap_8 FILLER_8_1722 ();
 sg13g2_decap_8 FILLER_8_1729 ();
 sg13g2_decap_8 FILLER_8_1736 ();
 sg13g2_decap_8 FILLER_8_1743 ();
 sg13g2_decap_8 FILLER_8_1750 ();
 sg13g2_decap_8 FILLER_8_1757 ();
 sg13g2_decap_8 FILLER_8_1764 ();
 sg13g2_decap_8 FILLER_8_1771 ();
 sg13g2_decap_8 FILLER_8_1778 ();
 sg13g2_decap_8 FILLER_8_1785 ();
 sg13g2_decap_8 FILLER_8_1792 ();
 sg13g2_decap_8 FILLER_8_1799 ();
 sg13g2_decap_8 FILLER_8_1806 ();
 sg13g2_decap_8 FILLER_8_1813 ();
 sg13g2_decap_8 FILLER_8_1820 ();
 sg13g2_decap_8 FILLER_8_1827 ();
 sg13g2_decap_8 FILLER_8_1834 ();
 sg13g2_decap_8 FILLER_8_1841 ();
 sg13g2_decap_8 FILLER_8_1848 ();
 sg13g2_decap_8 FILLER_8_1855 ();
 sg13g2_decap_8 FILLER_8_1862 ();
 sg13g2_decap_8 FILLER_8_1869 ();
 sg13g2_decap_8 FILLER_8_1876 ();
 sg13g2_decap_8 FILLER_8_1883 ();
 sg13g2_decap_8 FILLER_8_1890 ();
 sg13g2_decap_8 FILLER_8_1897 ();
 sg13g2_decap_8 FILLER_8_1904 ();
 sg13g2_decap_8 FILLER_8_1911 ();
 sg13g2_decap_8 FILLER_8_1918 ();
 sg13g2_decap_8 FILLER_8_1925 ();
 sg13g2_decap_8 FILLER_8_1932 ();
 sg13g2_decap_8 FILLER_8_1939 ();
 sg13g2_decap_8 FILLER_8_1946 ();
 sg13g2_decap_8 FILLER_8_1953 ();
 sg13g2_decap_8 FILLER_8_1960 ();
 sg13g2_decap_8 FILLER_8_1967 ();
 sg13g2_decap_8 FILLER_8_1974 ();
 sg13g2_decap_8 FILLER_8_1981 ();
 sg13g2_decap_8 FILLER_8_1988 ();
 sg13g2_decap_8 FILLER_8_1995 ();
 sg13g2_decap_8 FILLER_8_2002 ();
 sg13g2_decap_8 FILLER_8_2009 ();
 sg13g2_decap_8 FILLER_8_2016 ();
 sg13g2_decap_8 FILLER_8_2023 ();
 sg13g2_decap_8 FILLER_8_2030 ();
 sg13g2_decap_8 FILLER_8_2037 ();
 sg13g2_decap_8 FILLER_8_2044 ();
 sg13g2_fill_2 FILLER_8_2051 ();
 sg13g2_fill_1 FILLER_8_2053 ();
 sg13g2_decap_8 FILLER_8_2075 ();
 sg13g2_decap_8 FILLER_8_2082 ();
 sg13g2_decap_8 FILLER_8_2089 ();
 sg13g2_decap_8 FILLER_8_2096 ();
 sg13g2_decap_8 FILLER_8_2103 ();
 sg13g2_decap_8 FILLER_8_2110 ();
 sg13g2_decap_8 FILLER_8_2117 ();
 sg13g2_decap_8 FILLER_8_2124 ();
 sg13g2_decap_8 FILLER_8_2131 ();
 sg13g2_decap_8 FILLER_8_2138 ();
 sg13g2_decap_8 FILLER_8_2145 ();
 sg13g2_decap_8 FILLER_8_2152 ();
 sg13g2_decap_8 FILLER_8_2159 ();
 sg13g2_decap_8 FILLER_8_2166 ();
 sg13g2_decap_8 FILLER_8_2173 ();
 sg13g2_decap_8 FILLER_8_2180 ();
 sg13g2_decap_8 FILLER_8_2187 ();
 sg13g2_decap_8 FILLER_8_2194 ();
 sg13g2_decap_8 FILLER_8_2201 ();
 sg13g2_decap_4 FILLER_8_2208 ();
 sg13g2_decap_8 FILLER_8_2233 ();
 sg13g2_decap_8 FILLER_8_2240 ();
 sg13g2_decap_8 FILLER_8_2247 ();
 sg13g2_decap_4 FILLER_8_2254 ();
 sg13g2_fill_2 FILLER_8_2258 ();
 sg13g2_decap_8 FILLER_8_2275 ();
 sg13g2_decap_8 FILLER_8_2282 ();
 sg13g2_decap_8 FILLER_8_2289 ();
 sg13g2_decap_8 FILLER_8_2296 ();
 sg13g2_decap_8 FILLER_8_2303 ();
 sg13g2_decap_8 FILLER_8_2310 ();
 sg13g2_decap_8 FILLER_8_2317 ();
 sg13g2_decap_8 FILLER_8_2324 ();
 sg13g2_decap_8 FILLER_8_2331 ();
 sg13g2_fill_1 FILLER_8_2338 ();
 sg13g2_decap_8 FILLER_8_2364 ();
 sg13g2_decap_8 FILLER_8_2371 ();
 sg13g2_fill_2 FILLER_8_2378 ();
 sg13g2_fill_1 FILLER_8_2380 ();
 sg13g2_decap_8 FILLER_8_2406 ();
 sg13g2_decap_8 FILLER_8_2413 ();
 sg13g2_fill_2 FILLER_8_2420 ();
 sg13g2_decap_8 FILLER_8_2447 ();
 sg13g2_decap_8 FILLER_8_2454 ();
 sg13g2_decap_8 FILLER_8_2461 ();
 sg13g2_decap_8 FILLER_8_2468 ();
 sg13g2_decap_8 FILLER_8_2475 ();
 sg13g2_decap_8 FILLER_8_2482 ();
 sg13g2_fill_1 FILLER_8_2489 ();
 sg13g2_decap_8 FILLER_8_2515 ();
 sg13g2_decap_8 FILLER_8_2522 ();
 sg13g2_decap_8 FILLER_8_2529 ();
 sg13g2_decap_4 FILLER_8_2536 ();
 sg13g2_fill_1 FILLER_8_2540 ();
 sg13g2_decap_8 FILLER_8_2570 ();
 sg13g2_decap_8 FILLER_8_2577 ();
 sg13g2_decap_4 FILLER_8_2584 ();
 sg13g2_fill_2 FILLER_8_2588 ();
 sg13g2_decap_8 FILLER_8_2596 ();
 sg13g2_decap_8 FILLER_8_2603 ();
 sg13g2_decap_8 FILLER_8_2610 ();
 sg13g2_decap_8 FILLER_8_2617 ();
 sg13g2_decap_8 FILLER_8_2624 ();
 sg13g2_fill_1 FILLER_8_2631 ();
 sg13g2_decap_8 FILLER_8_2645 ();
 sg13g2_fill_2 FILLER_8_2652 ();
 sg13g2_decap_8 FILLER_8_2673 ();
 sg13g2_decap_4 FILLER_8_2680 ();
 sg13g2_decap_8 FILLER_8_2687 ();
 sg13g2_decap_4 FILLER_8_2694 ();
 sg13g2_fill_2 FILLER_8_2698 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_4 FILLER_9_826 ();
 sg13g2_fill_1 FILLER_9_830 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_decap_8 FILLER_9_863 ();
 sg13g2_decap_8 FILLER_9_870 ();
 sg13g2_decap_8 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_9_884 ();
 sg13g2_decap_8 FILLER_9_891 ();
 sg13g2_decap_8 FILLER_9_898 ();
 sg13g2_decap_8 FILLER_9_905 ();
 sg13g2_decap_8 FILLER_9_912 ();
 sg13g2_decap_8 FILLER_9_919 ();
 sg13g2_decap_8 FILLER_9_926 ();
 sg13g2_decap_8 FILLER_9_933 ();
 sg13g2_decap_8 FILLER_9_940 ();
 sg13g2_decap_8 FILLER_9_947 ();
 sg13g2_decap_8 FILLER_9_954 ();
 sg13g2_decap_8 FILLER_9_961 ();
 sg13g2_decap_8 FILLER_9_968 ();
 sg13g2_decap_8 FILLER_9_975 ();
 sg13g2_decap_8 FILLER_9_982 ();
 sg13g2_decap_8 FILLER_9_989 ();
 sg13g2_decap_8 FILLER_9_996 ();
 sg13g2_decap_8 FILLER_9_1003 ();
 sg13g2_decap_8 FILLER_9_1010 ();
 sg13g2_decap_8 FILLER_9_1017 ();
 sg13g2_decap_8 FILLER_9_1024 ();
 sg13g2_decap_8 FILLER_9_1031 ();
 sg13g2_decap_8 FILLER_9_1038 ();
 sg13g2_decap_8 FILLER_9_1045 ();
 sg13g2_decap_8 FILLER_9_1052 ();
 sg13g2_decap_8 FILLER_9_1059 ();
 sg13g2_decap_8 FILLER_9_1066 ();
 sg13g2_decap_8 FILLER_9_1073 ();
 sg13g2_decap_8 FILLER_9_1080 ();
 sg13g2_decap_8 FILLER_9_1087 ();
 sg13g2_decap_8 FILLER_9_1094 ();
 sg13g2_decap_8 FILLER_9_1101 ();
 sg13g2_decap_8 FILLER_9_1108 ();
 sg13g2_decap_8 FILLER_9_1115 ();
 sg13g2_decap_8 FILLER_9_1122 ();
 sg13g2_fill_2 FILLER_9_1129 ();
 sg13g2_decap_8 FILLER_9_1156 ();
 sg13g2_decap_8 FILLER_9_1163 ();
 sg13g2_fill_2 FILLER_9_1170 ();
 sg13g2_fill_1 FILLER_9_1172 ();
 sg13g2_decap_8 FILLER_9_1194 ();
 sg13g2_decap_8 FILLER_9_1201 ();
 sg13g2_decap_8 FILLER_9_1208 ();
 sg13g2_decap_8 FILLER_9_1215 ();
 sg13g2_decap_8 FILLER_9_1222 ();
 sg13g2_decap_8 FILLER_9_1229 ();
 sg13g2_decap_8 FILLER_9_1236 ();
 sg13g2_decap_8 FILLER_9_1243 ();
 sg13g2_fill_2 FILLER_9_1250 ();
 sg13g2_decap_8 FILLER_9_1277 ();
 sg13g2_fill_2 FILLER_9_1284 ();
 sg13g2_fill_1 FILLER_9_1286 ();
 sg13g2_decap_8 FILLER_9_1292 ();
 sg13g2_fill_2 FILLER_9_1299 ();
 sg13g2_decap_8 FILLER_9_1326 ();
 sg13g2_decap_8 FILLER_9_1333 ();
 sg13g2_decap_8 FILLER_9_1340 ();
 sg13g2_decap_8 FILLER_9_1347 ();
 sg13g2_decap_8 FILLER_9_1354 ();
 sg13g2_decap_8 FILLER_9_1361 ();
 sg13g2_decap_8 FILLER_9_1368 ();
 sg13g2_decap_8 FILLER_9_1375 ();
 sg13g2_decap_8 FILLER_9_1382 ();
 sg13g2_decap_8 FILLER_9_1389 ();
 sg13g2_decap_8 FILLER_9_1396 ();
 sg13g2_decap_8 FILLER_9_1403 ();
 sg13g2_decap_8 FILLER_9_1410 ();
 sg13g2_decap_8 FILLER_9_1417 ();
 sg13g2_decap_8 FILLER_9_1424 ();
 sg13g2_decap_8 FILLER_9_1431 ();
 sg13g2_decap_8 FILLER_9_1438 ();
 sg13g2_decap_8 FILLER_9_1445 ();
 sg13g2_decap_8 FILLER_9_1452 ();
 sg13g2_decap_4 FILLER_9_1459 ();
 sg13g2_decap_8 FILLER_9_1466 ();
 sg13g2_decap_8 FILLER_9_1473 ();
 sg13g2_decap_8 FILLER_9_1480 ();
 sg13g2_decap_8 FILLER_9_1487 ();
 sg13g2_decap_8 FILLER_9_1494 ();
 sg13g2_fill_1 FILLER_9_1501 ();
 sg13g2_decap_8 FILLER_9_1505 ();
 sg13g2_decap_8 FILLER_9_1512 ();
 sg13g2_decap_8 FILLER_9_1519 ();
 sg13g2_decap_8 FILLER_9_1526 ();
 sg13g2_decap_8 FILLER_9_1533 ();
 sg13g2_decap_8 FILLER_9_1540 ();
 sg13g2_decap_8 FILLER_9_1547 ();
 sg13g2_decap_8 FILLER_9_1554 ();
 sg13g2_decap_8 FILLER_9_1561 ();
 sg13g2_decap_8 FILLER_9_1568 ();
 sg13g2_decap_8 FILLER_9_1575 ();
 sg13g2_decap_8 FILLER_9_1582 ();
 sg13g2_decap_8 FILLER_9_1589 ();
 sg13g2_decap_8 FILLER_9_1596 ();
 sg13g2_decap_8 FILLER_9_1603 ();
 sg13g2_decap_8 FILLER_9_1610 ();
 sg13g2_decap_8 FILLER_9_1617 ();
 sg13g2_decap_8 FILLER_9_1624 ();
 sg13g2_decap_8 FILLER_9_1631 ();
 sg13g2_decap_8 FILLER_9_1638 ();
 sg13g2_decap_8 FILLER_9_1645 ();
 sg13g2_decap_8 FILLER_9_1652 ();
 sg13g2_decap_8 FILLER_9_1659 ();
 sg13g2_decap_8 FILLER_9_1666 ();
 sg13g2_decap_8 FILLER_9_1673 ();
 sg13g2_decap_8 FILLER_9_1680 ();
 sg13g2_decap_8 FILLER_9_1687 ();
 sg13g2_decap_8 FILLER_9_1694 ();
 sg13g2_decap_8 FILLER_9_1701 ();
 sg13g2_decap_8 FILLER_9_1708 ();
 sg13g2_decap_8 FILLER_9_1715 ();
 sg13g2_decap_8 FILLER_9_1722 ();
 sg13g2_decap_8 FILLER_9_1729 ();
 sg13g2_decap_8 FILLER_9_1736 ();
 sg13g2_decap_8 FILLER_9_1743 ();
 sg13g2_decap_8 FILLER_9_1750 ();
 sg13g2_decap_8 FILLER_9_1757 ();
 sg13g2_decap_8 FILLER_9_1764 ();
 sg13g2_decap_8 FILLER_9_1771 ();
 sg13g2_decap_8 FILLER_9_1778 ();
 sg13g2_decap_8 FILLER_9_1785 ();
 sg13g2_decap_8 FILLER_9_1792 ();
 sg13g2_decap_8 FILLER_9_1799 ();
 sg13g2_decap_8 FILLER_9_1806 ();
 sg13g2_decap_8 FILLER_9_1813 ();
 sg13g2_decap_8 FILLER_9_1820 ();
 sg13g2_decap_8 FILLER_9_1827 ();
 sg13g2_decap_8 FILLER_9_1834 ();
 sg13g2_decap_8 FILLER_9_1841 ();
 sg13g2_decap_8 FILLER_9_1848 ();
 sg13g2_decap_8 FILLER_9_1855 ();
 sg13g2_decap_8 FILLER_9_1862 ();
 sg13g2_decap_8 FILLER_9_1869 ();
 sg13g2_decap_8 FILLER_9_1876 ();
 sg13g2_decap_8 FILLER_9_1883 ();
 sg13g2_decap_8 FILLER_9_1890 ();
 sg13g2_decap_8 FILLER_9_1897 ();
 sg13g2_decap_8 FILLER_9_1904 ();
 sg13g2_decap_8 FILLER_9_1911 ();
 sg13g2_decap_8 FILLER_9_1918 ();
 sg13g2_decap_8 FILLER_9_1925 ();
 sg13g2_decap_4 FILLER_9_1932 ();
 sg13g2_fill_2 FILLER_9_1936 ();
 sg13g2_decap_8 FILLER_9_1943 ();
 sg13g2_decap_8 FILLER_9_1950 ();
 sg13g2_decap_8 FILLER_9_1957 ();
 sg13g2_decap_8 FILLER_9_1964 ();
 sg13g2_decap_8 FILLER_9_1971 ();
 sg13g2_decap_8 FILLER_9_1978 ();
 sg13g2_decap_8 FILLER_9_1985 ();
 sg13g2_decap_8 FILLER_9_1992 ();
 sg13g2_decap_8 FILLER_9_1999 ();
 sg13g2_decap_8 FILLER_9_2006 ();
 sg13g2_decap_8 FILLER_9_2013 ();
 sg13g2_decap_8 FILLER_9_2020 ();
 sg13g2_decap_8 FILLER_9_2027 ();
 sg13g2_decap_8 FILLER_9_2034 ();
 sg13g2_decap_8 FILLER_9_2041 ();
 sg13g2_decap_4 FILLER_9_2048 ();
 sg13g2_fill_1 FILLER_9_2052 ();
 sg13g2_decap_8 FILLER_9_2078 ();
 sg13g2_decap_8 FILLER_9_2085 ();
 sg13g2_decap_8 FILLER_9_2092 ();
 sg13g2_decap_8 FILLER_9_2099 ();
 sg13g2_decap_4 FILLER_9_2106 ();
 sg13g2_fill_1 FILLER_9_2110 ();
 sg13g2_decap_8 FILLER_9_2114 ();
 sg13g2_decap_8 FILLER_9_2121 ();
 sg13g2_decap_8 FILLER_9_2128 ();
 sg13g2_decap_8 FILLER_9_2135 ();
 sg13g2_decap_8 FILLER_9_2142 ();
 sg13g2_decap_8 FILLER_9_2149 ();
 sg13g2_decap_8 FILLER_9_2156 ();
 sg13g2_decap_8 FILLER_9_2163 ();
 sg13g2_fill_2 FILLER_9_2170 ();
 sg13g2_fill_1 FILLER_9_2172 ();
 sg13g2_decap_8 FILLER_9_2194 ();
 sg13g2_decap_8 FILLER_9_2201 ();
 sg13g2_decap_4 FILLER_9_2208 ();
 sg13g2_fill_1 FILLER_9_2212 ();
 sg13g2_decap_8 FILLER_9_2238 ();
 sg13g2_decap_8 FILLER_9_2245 ();
 sg13g2_decap_8 FILLER_9_2252 ();
 sg13g2_decap_8 FILLER_9_2259 ();
 sg13g2_decap_8 FILLER_9_2266 ();
 sg13g2_decap_8 FILLER_9_2273 ();
 sg13g2_decap_8 FILLER_9_2280 ();
 sg13g2_decap_8 FILLER_9_2287 ();
 sg13g2_decap_4 FILLER_9_2294 ();
 sg13g2_decap_8 FILLER_9_2313 ();
 sg13g2_fill_2 FILLER_9_2320 ();
 sg13g2_fill_1 FILLER_9_2322 ();
 sg13g2_decap_8 FILLER_9_2338 ();
 sg13g2_decap_8 FILLER_9_2345 ();
 sg13g2_decap_8 FILLER_9_2352 ();
 sg13g2_decap_8 FILLER_9_2359 ();
 sg13g2_decap_8 FILLER_9_2366 ();
 sg13g2_decap_8 FILLER_9_2373 ();
 sg13g2_decap_8 FILLER_9_2380 ();
 sg13g2_decap_8 FILLER_9_2387 ();
 sg13g2_decap_8 FILLER_9_2394 ();
 sg13g2_decap_8 FILLER_9_2401 ();
 sg13g2_decap_8 FILLER_9_2408 ();
 sg13g2_decap_8 FILLER_9_2415 ();
 sg13g2_decap_8 FILLER_9_2422 ();
 sg13g2_decap_8 FILLER_9_2429 ();
 sg13g2_decap_8 FILLER_9_2436 ();
 sg13g2_decap_8 FILLER_9_2443 ();
 sg13g2_decap_8 FILLER_9_2450 ();
 sg13g2_decap_8 FILLER_9_2457 ();
 sg13g2_decap_8 FILLER_9_2464 ();
 sg13g2_decap_8 FILLER_9_2471 ();
 sg13g2_decap_8 FILLER_9_2478 ();
 sg13g2_decap_8 FILLER_9_2485 ();
 sg13g2_decap_8 FILLER_9_2492 ();
 sg13g2_fill_1 FILLER_9_2499 ();
 sg13g2_decap_8 FILLER_9_2505 ();
 sg13g2_decap_8 FILLER_9_2512 ();
 sg13g2_decap_8 FILLER_9_2519 ();
 sg13g2_decap_4 FILLER_9_2526 ();
 sg13g2_fill_1 FILLER_9_2530 ();
 sg13g2_decap_8 FILLER_9_2540 ();
 sg13g2_decap_8 FILLER_9_2547 ();
 sg13g2_decap_4 FILLER_9_2554 ();
 sg13g2_decap_8 FILLER_9_2561 ();
 sg13g2_decap_8 FILLER_9_2568 ();
 sg13g2_decap_8 FILLER_9_2575 ();
 sg13g2_fill_2 FILLER_9_2582 ();
 sg13g2_fill_1 FILLER_9_2584 ();
 sg13g2_decap_8 FILLER_9_2601 ();
 sg13g2_fill_2 FILLER_9_2608 ();
 sg13g2_decap_4 FILLER_9_2632 ();
 sg13g2_fill_1 FILLER_9_2636 ();
 sg13g2_fill_2 FILLER_9_2643 ();
 sg13g2_decap_8 FILLER_9_2648 ();
 sg13g2_decap_8 FILLER_9_2655 ();
 sg13g2_decap_8 FILLER_9_2662 ();
 sg13g2_decap_8 FILLER_9_2669 ();
 sg13g2_decap_8 FILLER_9_2676 ();
 sg13g2_fill_1 FILLER_9_2683 ();
 sg13g2_decap_8 FILLER_9_2687 ();
 sg13g2_decap_4 FILLER_9_2694 ();
 sg13g2_fill_2 FILLER_9_2698 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_4 FILLER_10_651 ();
 sg13g2_fill_2 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_660 ();
 sg13g2_decap_8 FILLER_10_667 ();
 sg13g2_decap_8 FILLER_10_674 ();
 sg13g2_fill_2 FILLER_10_681 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_872 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_decap_4 FILLER_10_886 ();
 sg13g2_decap_8 FILLER_10_915 ();
 sg13g2_decap_8 FILLER_10_922 ();
 sg13g2_decap_8 FILLER_10_929 ();
 sg13g2_decap_8 FILLER_10_936 ();
 sg13g2_decap_8 FILLER_10_943 ();
 sg13g2_decap_8 FILLER_10_950 ();
 sg13g2_decap_8 FILLER_10_957 ();
 sg13g2_fill_1 FILLER_10_964 ();
 sg13g2_decap_8 FILLER_10_975 ();
 sg13g2_decap_8 FILLER_10_982 ();
 sg13g2_decap_8 FILLER_10_989 ();
 sg13g2_decap_8 FILLER_10_996 ();
 sg13g2_decap_8 FILLER_10_1003 ();
 sg13g2_decap_8 FILLER_10_1010 ();
 sg13g2_fill_1 FILLER_10_1017 ();
 sg13g2_decap_8 FILLER_10_1039 ();
 sg13g2_decap_8 FILLER_10_1046 ();
 sg13g2_decap_8 FILLER_10_1053 ();
 sg13g2_decap_8 FILLER_10_1081 ();
 sg13g2_decap_8 FILLER_10_1088 ();
 sg13g2_decap_4 FILLER_10_1095 ();
 sg13g2_decap_8 FILLER_10_1120 ();
 sg13g2_decap_8 FILLER_10_1127 ();
 sg13g2_decap_8 FILLER_10_1134 ();
 sg13g2_decap_8 FILLER_10_1141 ();
 sg13g2_decap_8 FILLER_10_1148 ();
 sg13g2_decap_8 FILLER_10_1155 ();
 sg13g2_decap_8 FILLER_10_1162 ();
 sg13g2_decap_8 FILLER_10_1169 ();
 sg13g2_decap_8 FILLER_10_1176 ();
 sg13g2_decap_8 FILLER_10_1183 ();
 sg13g2_decap_8 FILLER_10_1190 ();
 sg13g2_decap_8 FILLER_10_1197 ();
 sg13g2_decap_8 FILLER_10_1204 ();
 sg13g2_decap_8 FILLER_10_1211 ();
 sg13g2_decap_8 FILLER_10_1218 ();
 sg13g2_decap_8 FILLER_10_1225 ();
 sg13g2_decap_8 FILLER_10_1232 ();
 sg13g2_decap_8 FILLER_10_1239 ();
 sg13g2_decap_8 FILLER_10_1246 ();
 sg13g2_decap_8 FILLER_10_1253 ();
 sg13g2_decap_8 FILLER_10_1260 ();
 sg13g2_decap_8 FILLER_10_1267 ();
 sg13g2_decap_8 FILLER_10_1274 ();
 sg13g2_decap_8 FILLER_10_1281 ();
 sg13g2_decap_8 FILLER_10_1288 ();
 sg13g2_decap_8 FILLER_10_1295 ();
 sg13g2_decap_8 FILLER_10_1302 ();
 sg13g2_decap_8 FILLER_10_1309 ();
 sg13g2_decap_8 FILLER_10_1316 ();
 sg13g2_decap_8 FILLER_10_1323 ();
 sg13g2_decap_8 FILLER_10_1330 ();
 sg13g2_decap_8 FILLER_10_1337 ();
 sg13g2_decap_8 FILLER_10_1344 ();
 sg13g2_decap_8 FILLER_10_1351 ();
 sg13g2_decap_8 FILLER_10_1358 ();
 sg13g2_decap_8 FILLER_10_1365 ();
 sg13g2_decap_8 FILLER_10_1372 ();
 sg13g2_decap_8 FILLER_10_1379 ();
 sg13g2_decap_8 FILLER_10_1386 ();
 sg13g2_decap_8 FILLER_10_1393 ();
 sg13g2_decap_8 FILLER_10_1400 ();
 sg13g2_decap_8 FILLER_10_1407 ();
 sg13g2_decap_8 FILLER_10_1414 ();
 sg13g2_decap_8 FILLER_10_1421 ();
 sg13g2_decap_8 FILLER_10_1428 ();
 sg13g2_decap_8 FILLER_10_1435 ();
 sg13g2_decap_8 FILLER_10_1442 ();
 sg13g2_decap_8 FILLER_10_1449 ();
 sg13g2_decap_8 FILLER_10_1456 ();
 sg13g2_decap_8 FILLER_10_1463 ();
 sg13g2_decap_8 FILLER_10_1470 ();
 sg13g2_decap_8 FILLER_10_1477 ();
 sg13g2_decap_8 FILLER_10_1484 ();
 sg13g2_decap_8 FILLER_10_1491 ();
 sg13g2_decap_8 FILLER_10_1498 ();
 sg13g2_decap_4 FILLER_10_1505 ();
 sg13g2_fill_1 FILLER_10_1509 ();
 sg13g2_decap_8 FILLER_10_1513 ();
 sg13g2_decap_4 FILLER_10_1520 ();
 sg13g2_fill_1 FILLER_10_1524 ();
 sg13g2_decap_8 FILLER_10_1528 ();
 sg13g2_decap_8 FILLER_10_1535 ();
 sg13g2_decap_8 FILLER_10_1542 ();
 sg13g2_decap_8 FILLER_10_1549 ();
 sg13g2_decap_8 FILLER_10_1556 ();
 sg13g2_decap_8 FILLER_10_1563 ();
 sg13g2_decap_8 FILLER_10_1570 ();
 sg13g2_decap_4 FILLER_10_1577 ();
 sg13g2_fill_1 FILLER_10_1581 ();
 sg13g2_decap_8 FILLER_10_1585 ();
 sg13g2_decap_8 FILLER_10_1592 ();
 sg13g2_decap_8 FILLER_10_1599 ();
 sg13g2_decap_8 FILLER_10_1606 ();
 sg13g2_decap_8 FILLER_10_1613 ();
 sg13g2_decap_8 FILLER_10_1620 ();
 sg13g2_decap_8 FILLER_10_1627 ();
 sg13g2_decap_8 FILLER_10_1634 ();
 sg13g2_decap_8 FILLER_10_1641 ();
 sg13g2_decap_8 FILLER_10_1648 ();
 sg13g2_decap_8 FILLER_10_1655 ();
 sg13g2_decap_8 FILLER_10_1662 ();
 sg13g2_decap_8 FILLER_10_1669 ();
 sg13g2_decap_8 FILLER_10_1676 ();
 sg13g2_decap_8 FILLER_10_1683 ();
 sg13g2_decap_8 FILLER_10_1690 ();
 sg13g2_decap_8 FILLER_10_1697 ();
 sg13g2_decap_8 FILLER_10_1704 ();
 sg13g2_decap_8 FILLER_10_1711 ();
 sg13g2_decap_8 FILLER_10_1718 ();
 sg13g2_decap_8 FILLER_10_1725 ();
 sg13g2_decap_8 FILLER_10_1732 ();
 sg13g2_decap_8 FILLER_10_1739 ();
 sg13g2_decap_8 FILLER_10_1746 ();
 sg13g2_decap_8 FILLER_10_1753 ();
 sg13g2_decap_8 FILLER_10_1760 ();
 sg13g2_decap_8 FILLER_10_1767 ();
 sg13g2_decap_8 FILLER_10_1774 ();
 sg13g2_decap_8 FILLER_10_1781 ();
 sg13g2_decap_8 FILLER_10_1788 ();
 sg13g2_decap_8 FILLER_10_1795 ();
 sg13g2_decap_8 FILLER_10_1802 ();
 sg13g2_decap_8 FILLER_10_1809 ();
 sg13g2_decap_8 FILLER_10_1816 ();
 sg13g2_decap_8 FILLER_10_1823 ();
 sg13g2_decap_8 FILLER_10_1830 ();
 sg13g2_decap_8 FILLER_10_1837 ();
 sg13g2_decap_8 FILLER_10_1844 ();
 sg13g2_decap_8 FILLER_10_1851 ();
 sg13g2_decap_8 FILLER_10_1858 ();
 sg13g2_decap_8 FILLER_10_1865 ();
 sg13g2_decap_8 FILLER_10_1872 ();
 sg13g2_decap_8 FILLER_10_1879 ();
 sg13g2_decap_8 FILLER_10_1886 ();
 sg13g2_decap_8 FILLER_10_1893 ();
 sg13g2_decap_8 FILLER_10_1900 ();
 sg13g2_decap_8 FILLER_10_1907 ();
 sg13g2_decap_8 FILLER_10_1914 ();
 sg13g2_decap_8 FILLER_10_1921 ();
 sg13g2_decap_8 FILLER_10_1949 ();
 sg13g2_decap_8 FILLER_10_1956 ();
 sg13g2_decap_8 FILLER_10_1963 ();
 sg13g2_fill_1 FILLER_10_1970 ();
 sg13g2_decap_8 FILLER_10_1992 ();
 sg13g2_decap_8 FILLER_10_1999 ();
 sg13g2_decap_8 FILLER_10_2006 ();
 sg13g2_decap_4 FILLER_10_2013 ();
 sg13g2_decap_8 FILLER_10_2038 ();
 sg13g2_decap_8 FILLER_10_2045 ();
 sg13g2_decap_8 FILLER_10_2052 ();
 sg13g2_decap_8 FILLER_10_2059 ();
 sg13g2_decap_8 FILLER_10_2066 ();
 sg13g2_decap_8 FILLER_10_2073 ();
 sg13g2_decap_8 FILLER_10_2080 ();
 sg13g2_decap_8 FILLER_10_2087 ();
 sg13g2_fill_2 FILLER_10_2094 ();
 sg13g2_fill_1 FILLER_10_2096 ();
 sg13g2_decap_8 FILLER_10_2118 ();
 sg13g2_decap_8 FILLER_10_2125 ();
 sg13g2_decap_8 FILLER_10_2132 ();
 sg13g2_decap_8 FILLER_10_2139 ();
 sg13g2_decap_8 FILLER_10_2146 ();
 sg13g2_decap_8 FILLER_10_2153 ();
 sg13g2_decap_8 FILLER_10_2160 ();
 sg13g2_fill_2 FILLER_10_2167 ();
 sg13g2_decap_8 FILLER_10_2194 ();
 sg13g2_decap_8 FILLER_10_2201 ();
 sg13g2_decap_8 FILLER_10_2208 ();
 sg13g2_decap_8 FILLER_10_2215 ();
 sg13g2_decap_8 FILLER_10_2222 ();
 sg13g2_decap_8 FILLER_10_2229 ();
 sg13g2_decap_8 FILLER_10_2236 ();
 sg13g2_decap_8 FILLER_10_2243 ();
 sg13g2_decap_8 FILLER_10_2250 ();
 sg13g2_decap_4 FILLER_10_2257 ();
 sg13g2_decap_8 FILLER_10_2276 ();
 sg13g2_decap_8 FILLER_10_2283 ();
 sg13g2_decap_8 FILLER_10_2290 ();
 sg13g2_fill_2 FILLER_10_2297 ();
 sg13g2_fill_1 FILLER_10_2299 ();
 sg13g2_decap_8 FILLER_10_2315 ();
 sg13g2_decap_8 FILLER_10_2322 ();
 sg13g2_decap_8 FILLER_10_2329 ();
 sg13g2_decap_8 FILLER_10_2336 ();
 sg13g2_decap_8 FILLER_10_2343 ();
 sg13g2_decap_8 FILLER_10_2350 ();
 sg13g2_decap_8 FILLER_10_2357 ();
 sg13g2_decap_8 FILLER_10_2364 ();
 sg13g2_decap_8 FILLER_10_2371 ();
 sg13g2_decap_8 FILLER_10_2378 ();
 sg13g2_fill_2 FILLER_10_2385 ();
 sg13g2_fill_1 FILLER_10_2387 ();
 sg13g2_decap_8 FILLER_10_2393 ();
 sg13g2_decap_8 FILLER_10_2400 ();
 sg13g2_decap_8 FILLER_10_2407 ();
 sg13g2_decap_8 FILLER_10_2414 ();
 sg13g2_decap_8 FILLER_10_2421 ();
 sg13g2_decap_4 FILLER_10_2453 ();
 sg13g2_fill_2 FILLER_10_2457 ();
 sg13g2_decap_8 FILLER_10_2484 ();
 sg13g2_decap_8 FILLER_10_2491 ();
 sg13g2_decap_8 FILLER_10_2498 ();
 sg13g2_decap_8 FILLER_10_2505 ();
 sg13g2_decap_8 FILLER_10_2512 ();
 sg13g2_decap_8 FILLER_10_2519 ();
 sg13g2_fill_2 FILLER_10_2526 ();
 sg13g2_decap_8 FILLER_10_2541 ();
 sg13g2_decap_8 FILLER_10_2548 ();
 sg13g2_decap_4 FILLER_10_2555 ();
 sg13g2_fill_2 FILLER_10_2559 ();
 sg13g2_decap_8 FILLER_10_2564 ();
 sg13g2_decap_8 FILLER_10_2571 ();
 sg13g2_decap_8 FILLER_10_2578 ();
 sg13g2_fill_2 FILLER_10_2585 ();
 sg13g2_fill_1 FILLER_10_2587 ();
 sg13g2_decap_8 FILLER_10_2591 ();
 sg13g2_decap_8 FILLER_10_2598 ();
 sg13g2_decap_8 FILLER_10_2605 ();
 sg13g2_decap_8 FILLER_10_2612 ();
 sg13g2_decap_8 FILLER_10_2619 ();
 sg13g2_decap_8 FILLER_10_2626 ();
 sg13g2_decap_8 FILLER_10_2633 ();
 sg13g2_decap_8 FILLER_10_2640 ();
 sg13g2_decap_8 FILLER_10_2647 ();
 sg13g2_decap_8 FILLER_10_2654 ();
 sg13g2_decap_8 FILLER_10_2661 ();
 sg13g2_decap_8 FILLER_10_2668 ();
 sg13g2_decap_8 FILLER_10_2675 ();
 sg13g2_decap_8 FILLER_10_2682 ();
 sg13g2_decap_8 FILLER_10_2689 ();
 sg13g2_decap_4 FILLER_10_2696 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_4 FILLER_11_546 ();
 sg13g2_fill_2 FILLER_11_550 ();
 sg13g2_decap_8 FILLER_11_573 ();
 sg13g2_decap_8 FILLER_11_580 ();
 sg13g2_decap_8 FILLER_11_587 ();
 sg13g2_fill_2 FILLER_11_594 ();
 sg13g2_fill_1 FILLER_11_596 ();
 sg13g2_fill_1 FILLER_11_618 ();
 sg13g2_decap_8 FILLER_11_640 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_decap_8 FILLER_11_654 ();
 sg13g2_decap_8 FILLER_11_661 ();
 sg13g2_decap_8 FILLER_11_668 ();
 sg13g2_decap_8 FILLER_11_675 ();
 sg13g2_decap_8 FILLER_11_682 ();
 sg13g2_decap_8 FILLER_11_689 ();
 sg13g2_decap_8 FILLER_11_696 ();
 sg13g2_decap_8 FILLER_11_703 ();
 sg13g2_decap_8 FILLER_11_710 ();
 sg13g2_decap_8 FILLER_11_717 ();
 sg13g2_decap_8 FILLER_11_724 ();
 sg13g2_decap_8 FILLER_11_731 ();
 sg13g2_decap_4 FILLER_11_738 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_fill_2 FILLER_11_851 ();
 sg13g2_fill_1 FILLER_11_853 ();
 sg13g2_decap_8 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_decap_8 FILLER_11_900 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_4 FILLER_11_921 ();
 sg13g2_fill_1 FILLER_11_925 ();
 sg13g2_decap_8 FILLER_11_951 ();
 sg13g2_decap_8 FILLER_11_958 ();
 sg13g2_decap_8 FILLER_11_965 ();
 sg13g2_decap_8 FILLER_11_972 ();
 sg13g2_decap_8 FILLER_11_979 ();
 sg13g2_decap_8 FILLER_11_986 ();
 sg13g2_decap_8 FILLER_11_993 ();
 sg13g2_decap_8 FILLER_11_1000 ();
 sg13g2_decap_4 FILLER_11_1007 ();
 sg13g2_decap_8 FILLER_11_1036 ();
 sg13g2_decap_8 FILLER_11_1043 ();
 sg13g2_decap_4 FILLER_11_1050 ();
 sg13g2_decap_8 FILLER_11_1079 ();
 sg13g2_decap_8 FILLER_11_1086 ();
 sg13g2_decap_4 FILLER_11_1093 ();
 sg13g2_decap_8 FILLER_11_1122 ();
 sg13g2_decap_8 FILLER_11_1129 ();
 sg13g2_decap_8 FILLER_11_1136 ();
 sg13g2_decap_8 FILLER_11_1143 ();
 sg13g2_decap_8 FILLER_11_1150 ();
 sg13g2_decap_8 FILLER_11_1157 ();
 sg13g2_decap_8 FILLER_11_1164 ();
 sg13g2_decap_8 FILLER_11_1171 ();
 sg13g2_decap_8 FILLER_11_1178 ();
 sg13g2_decap_8 FILLER_11_1185 ();
 sg13g2_decap_8 FILLER_11_1192 ();
 sg13g2_decap_8 FILLER_11_1220 ();
 sg13g2_decap_8 FILLER_11_1227 ();
 sg13g2_decap_4 FILLER_11_1234 ();
 sg13g2_fill_2 FILLER_11_1238 ();
 sg13g2_decap_8 FILLER_11_1261 ();
 sg13g2_decap_8 FILLER_11_1268 ();
 sg13g2_decap_8 FILLER_11_1275 ();
 sg13g2_decap_8 FILLER_11_1282 ();
 sg13g2_decap_8 FILLER_11_1289 ();
 sg13g2_decap_8 FILLER_11_1296 ();
 sg13g2_decap_8 FILLER_11_1303 ();
 sg13g2_decap_8 FILLER_11_1310 ();
 sg13g2_decap_8 FILLER_11_1317 ();
 sg13g2_decap_8 FILLER_11_1324 ();
 sg13g2_decap_8 FILLER_11_1331 ();
 sg13g2_decap_8 FILLER_11_1338 ();
 sg13g2_decap_8 FILLER_11_1345 ();
 sg13g2_decap_8 FILLER_11_1352 ();
 sg13g2_decap_8 FILLER_11_1359 ();
 sg13g2_decap_8 FILLER_11_1366 ();
 sg13g2_decap_8 FILLER_11_1373 ();
 sg13g2_decap_8 FILLER_11_1380 ();
 sg13g2_decap_8 FILLER_11_1387 ();
 sg13g2_decap_8 FILLER_11_1394 ();
 sg13g2_decap_8 FILLER_11_1401 ();
 sg13g2_decap_8 FILLER_11_1408 ();
 sg13g2_decap_8 FILLER_11_1415 ();
 sg13g2_decap_8 FILLER_11_1422 ();
 sg13g2_decap_8 FILLER_11_1429 ();
 sg13g2_decap_8 FILLER_11_1436 ();
 sg13g2_decap_8 FILLER_11_1443 ();
 sg13g2_decap_8 FILLER_11_1450 ();
 sg13g2_decap_8 FILLER_11_1457 ();
 sg13g2_decap_8 FILLER_11_1464 ();
 sg13g2_decap_8 FILLER_11_1471 ();
 sg13g2_decap_8 FILLER_11_1478 ();
 sg13g2_decap_8 FILLER_11_1485 ();
 sg13g2_decap_8 FILLER_11_1492 ();
 sg13g2_decap_8 FILLER_11_1499 ();
 sg13g2_decap_8 FILLER_11_1506 ();
 sg13g2_decap_8 FILLER_11_1513 ();
 sg13g2_decap_8 FILLER_11_1520 ();
 sg13g2_decap_8 FILLER_11_1527 ();
 sg13g2_decap_8 FILLER_11_1534 ();
 sg13g2_decap_8 FILLER_11_1541 ();
 sg13g2_decap_8 FILLER_11_1548 ();
 sg13g2_fill_2 FILLER_11_1555 ();
 sg13g2_decap_8 FILLER_11_1560 ();
 sg13g2_decap_8 FILLER_11_1567 ();
 sg13g2_decap_8 FILLER_11_1574 ();
 sg13g2_decap_8 FILLER_11_1581 ();
 sg13g2_decap_8 FILLER_11_1588 ();
 sg13g2_decap_8 FILLER_11_1595 ();
 sg13g2_decap_8 FILLER_11_1602 ();
 sg13g2_decap_8 FILLER_11_1609 ();
 sg13g2_decap_8 FILLER_11_1616 ();
 sg13g2_decap_8 FILLER_11_1623 ();
 sg13g2_decap_8 FILLER_11_1630 ();
 sg13g2_decap_8 FILLER_11_1637 ();
 sg13g2_decap_8 FILLER_11_1644 ();
 sg13g2_decap_8 FILLER_11_1651 ();
 sg13g2_decap_8 FILLER_11_1658 ();
 sg13g2_decap_8 FILLER_11_1665 ();
 sg13g2_decap_8 FILLER_11_1672 ();
 sg13g2_decap_8 FILLER_11_1679 ();
 sg13g2_decap_8 FILLER_11_1686 ();
 sg13g2_decap_8 FILLER_11_1693 ();
 sg13g2_decap_8 FILLER_11_1700 ();
 sg13g2_decap_8 FILLER_11_1707 ();
 sg13g2_decap_8 FILLER_11_1714 ();
 sg13g2_decap_8 FILLER_11_1721 ();
 sg13g2_decap_8 FILLER_11_1728 ();
 sg13g2_decap_8 FILLER_11_1735 ();
 sg13g2_decap_8 FILLER_11_1742 ();
 sg13g2_decap_8 FILLER_11_1749 ();
 sg13g2_decap_8 FILLER_11_1756 ();
 sg13g2_decap_8 FILLER_11_1763 ();
 sg13g2_decap_8 FILLER_11_1770 ();
 sg13g2_decap_8 FILLER_11_1777 ();
 sg13g2_decap_8 FILLER_11_1784 ();
 sg13g2_decap_8 FILLER_11_1791 ();
 sg13g2_decap_8 FILLER_11_1798 ();
 sg13g2_decap_8 FILLER_11_1805 ();
 sg13g2_decap_8 FILLER_11_1812 ();
 sg13g2_decap_8 FILLER_11_1819 ();
 sg13g2_decap_8 FILLER_11_1826 ();
 sg13g2_decap_8 FILLER_11_1833 ();
 sg13g2_decap_8 FILLER_11_1840 ();
 sg13g2_decap_8 FILLER_11_1847 ();
 sg13g2_decap_8 FILLER_11_1854 ();
 sg13g2_decap_8 FILLER_11_1861 ();
 sg13g2_decap_8 FILLER_11_1868 ();
 sg13g2_decap_8 FILLER_11_1875 ();
 sg13g2_decap_8 FILLER_11_1882 ();
 sg13g2_decap_8 FILLER_11_1889 ();
 sg13g2_decap_8 FILLER_11_1896 ();
 sg13g2_decap_8 FILLER_11_1903 ();
 sg13g2_decap_8 FILLER_11_1910 ();
 sg13g2_decap_8 FILLER_11_1917 ();
 sg13g2_decap_8 FILLER_11_1949 ();
 sg13g2_decap_8 FILLER_11_1956 ();
 sg13g2_decap_8 FILLER_11_1963 ();
 sg13g2_decap_8 FILLER_11_1995 ();
 sg13g2_decap_8 FILLER_11_2002 ();
 sg13g2_decap_4 FILLER_11_2009 ();
 sg13g2_decap_8 FILLER_11_2038 ();
 sg13g2_decap_8 FILLER_11_2045 ();
 sg13g2_decap_8 FILLER_11_2052 ();
 sg13g2_decap_8 FILLER_11_2059 ();
 sg13g2_decap_8 FILLER_11_2066 ();
 sg13g2_decap_8 FILLER_11_2073 ();
 sg13g2_decap_8 FILLER_11_2080 ();
 sg13g2_decap_8 FILLER_11_2087 ();
 sg13g2_fill_1 FILLER_11_2094 ();
 sg13g2_decap_8 FILLER_11_2120 ();
 sg13g2_decap_8 FILLER_11_2127 ();
 sg13g2_decap_4 FILLER_11_2134 ();
 sg13g2_decap_8 FILLER_11_2159 ();
 sg13g2_decap_8 FILLER_11_2166 ();
 sg13g2_decap_8 FILLER_11_2173 ();
 sg13g2_decap_8 FILLER_11_2180 ();
 sg13g2_decap_8 FILLER_11_2187 ();
 sg13g2_decap_8 FILLER_11_2194 ();
 sg13g2_decap_8 FILLER_11_2204 ();
 sg13g2_decap_8 FILLER_11_2211 ();
 sg13g2_decap_8 FILLER_11_2218 ();
 sg13g2_decap_8 FILLER_11_2225 ();
 sg13g2_decap_8 FILLER_11_2232 ();
 sg13g2_decap_8 FILLER_11_2239 ();
 sg13g2_decap_8 FILLER_11_2246 ();
 sg13g2_decap_8 FILLER_11_2253 ();
 sg13g2_fill_1 FILLER_11_2260 ();
 sg13g2_decap_8 FILLER_11_2276 ();
 sg13g2_decap_8 FILLER_11_2283 ();
 sg13g2_decap_8 FILLER_11_2290 ();
 sg13g2_fill_2 FILLER_11_2297 ();
 sg13g2_decap_8 FILLER_11_2314 ();
 sg13g2_decap_8 FILLER_11_2321 ();
 sg13g2_decap_8 FILLER_11_2328 ();
 sg13g2_decap_8 FILLER_11_2335 ();
 sg13g2_decap_4 FILLER_11_2342 ();
 sg13g2_decap_8 FILLER_11_2371 ();
 sg13g2_decap_8 FILLER_11_2403 ();
 sg13g2_decap_8 FILLER_11_2410 ();
 sg13g2_decap_8 FILLER_11_2417 ();
 sg13g2_decap_8 FILLER_11_2424 ();
 sg13g2_decap_8 FILLER_11_2431 ();
 sg13g2_fill_2 FILLER_11_2438 ();
 sg13g2_decap_8 FILLER_11_2445 ();
 sg13g2_decap_8 FILLER_11_2452 ();
 sg13g2_decap_8 FILLER_11_2459 ();
 sg13g2_decap_4 FILLER_11_2466 ();
 sg13g2_decap_8 FILLER_11_2475 ();
 sg13g2_decap_8 FILLER_11_2482 ();
 sg13g2_decap_8 FILLER_11_2489 ();
 sg13g2_decap_8 FILLER_11_2496 ();
 sg13g2_decap_4 FILLER_11_2503 ();
 sg13g2_fill_1 FILLER_11_2507 ();
 sg13g2_decap_8 FILLER_11_2513 ();
 sg13g2_decap_8 FILLER_11_2520 ();
 sg13g2_decap_8 FILLER_11_2527 ();
 sg13g2_decap_8 FILLER_11_2534 ();
 sg13g2_decap_8 FILLER_11_2541 ();
 sg13g2_decap_8 FILLER_11_2548 ();
 sg13g2_decap_8 FILLER_11_2561 ();
 sg13g2_decap_8 FILLER_11_2568 ();
 sg13g2_decap_8 FILLER_11_2575 ();
 sg13g2_decap_8 FILLER_11_2582 ();
 sg13g2_decap_8 FILLER_11_2589 ();
 sg13g2_fill_1 FILLER_11_2596 ();
 sg13g2_decap_8 FILLER_11_2600 ();
 sg13g2_decap_8 FILLER_11_2607 ();
 sg13g2_decap_8 FILLER_11_2614 ();
 sg13g2_fill_1 FILLER_11_2621 ();
 sg13g2_fill_2 FILLER_11_2628 ();
 sg13g2_decap_8 FILLER_11_2633 ();
 sg13g2_decap_8 FILLER_11_2640 ();
 sg13g2_decap_8 FILLER_11_2647 ();
 sg13g2_decap_8 FILLER_11_2654 ();
 sg13g2_decap_8 FILLER_11_2661 ();
 sg13g2_decap_8 FILLER_11_2668 ();
 sg13g2_decap_4 FILLER_11_2675 ();
 sg13g2_fill_1 FILLER_11_2679 ();
 sg13g2_decap_8 FILLER_11_2691 ();
 sg13g2_fill_2 FILLER_11_2698 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_fill_2 FILLER_12_686 ();
 sg13g2_fill_1 FILLER_12_688 ();
 sg13g2_decap_8 FILLER_12_710 ();
 sg13g2_decap_8 FILLER_12_717 ();
 sg13g2_decap_8 FILLER_12_724 ();
 sg13g2_decap_8 FILLER_12_731 ();
 sg13g2_decap_8 FILLER_12_738 ();
 sg13g2_decap_8 FILLER_12_745 ();
 sg13g2_decap_8 FILLER_12_752 ();
 sg13g2_decap_8 FILLER_12_759 ();
 sg13g2_decap_8 FILLER_12_766 ();
 sg13g2_decap_8 FILLER_12_773 ();
 sg13g2_decap_8 FILLER_12_780 ();
 sg13g2_decap_8 FILLER_12_787 ();
 sg13g2_decap_8 FILLER_12_794 ();
 sg13g2_decap_8 FILLER_12_801 ();
 sg13g2_decap_8 FILLER_12_808 ();
 sg13g2_decap_8 FILLER_12_815 ();
 sg13g2_decap_8 FILLER_12_822 ();
 sg13g2_fill_2 FILLER_12_829 ();
 sg13g2_decap_8 FILLER_12_856 ();
 sg13g2_decap_8 FILLER_12_863 ();
 sg13g2_decap_8 FILLER_12_870 ();
 sg13g2_decap_8 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_12_884 ();
 sg13g2_decap_8 FILLER_12_891 ();
 sg13g2_decap_8 FILLER_12_898 ();
 sg13g2_decap_8 FILLER_12_905 ();
 sg13g2_decap_8 FILLER_12_912 ();
 sg13g2_decap_8 FILLER_12_919 ();
 sg13g2_decap_8 FILLER_12_926 ();
 sg13g2_decap_8 FILLER_12_933 ();
 sg13g2_decap_8 FILLER_12_940 ();
 sg13g2_decap_8 FILLER_12_947 ();
 sg13g2_decap_8 FILLER_12_954 ();
 sg13g2_decap_8 FILLER_12_961 ();
 sg13g2_decap_8 FILLER_12_968 ();
 sg13g2_decap_8 FILLER_12_975 ();
 sg13g2_decap_8 FILLER_12_982 ();
 sg13g2_decap_8 FILLER_12_989 ();
 sg13g2_decap_8 FILLER_12_996 ();
 sg13g2_decap_8 FILLER_12_1003 ();
 sg13g2_decap_8 FILLER_12_1010 ();
 sg13g2_decap_8 FILLER_12_1017 ();
 sg13g2_decap_8 FILLER_12_1024 ();
 sg13g2_decap_8 FILLER_12_1031 ();
 sg13g2_decap_8 FILLER_12_1038 ();
 sg13g2_decap_8 FILLER_12_1045 ();
 sg13g2_decap_8 FILLER_12_1052 ();
 sg13g2_decap_8 FILLER_12_1059 ();
 sg13g2_decap_8 FILLER_12_1066 ();
 sg13g2_decap_8 FILLER_12_1073 ();
 sg13g2_decap_8 FILLER_12_1080 ();
 sg13g2_decap_8 FILLER_12_1087 ();
 sg13g2_decap_8 FILLER_12_1094 ();
 sg13g2_decap_8 FILLER_12_1101 ();
 sg13g2_decap_8 FILLER_12_1108 ();
 sg13g2_decap_8 FILLER_12_1115 ();
 sg13g2_decap_8 FILLER_12_1122 ();
 sg13g2_decap_8 FILLER_12_1129 ();
 sg13g2_decap_8 FILLER_12_1136 ();
 sg13g2_decap_8 FILLER_12_1143 ();
 sg13g2_decap_8 FILLER_12_1150 ();
 sg13g2_decap_8 FILLER_12_1157 ();
 sg13g2_decap_8 FILLER_12_1164 ();
 sg13g2_decap_8 FILLER_12_1171 ();
 sg13g2_decap_8 FILLER_12_1178 ();
 sg13g2_decap_8 FILLER_12_1185 ();
 sg13g2_decap_4 FILLER_12_1192 ();
 sg13g2_fill_1 FILLER_12_1196 ();
 sg13g2_decap_8 FILLER_12_1222 ();
 sg13g2_decap_8 FILLER_12_1229 ();
 sg13g2_fill_2 FILLER_12_1236 ();
 sg13g2_decap_8 FILLER_12_1263 ();
 sg13g2_decap_8 FILLER_12_1270 ();
 sg13g2_decap_8 FILLER_12_1277 ();
 sg13g2_fill_2 FILLER_12_1284 ();
 sg13g2_fill_1 FILLER_12_1286 ();
 sg13g2_decap_8 FILLER_12_1308 ();
 sg13g2_decap_4 FILLER_12_1315 ();
 sg13g2_fill_2 FILLER_12_1324 ();
 sg13g2_fill_1 FILLER_12_1326 ();
 sg13g2_decap_8 FILLER_12_1337 ();
 sg13g2_decap_8 FILLER_12_1344 ();
 sg13g2_decap_8 FILLER_12_1351 ();
 sg13g2_decap_8 FILLER_12_1358 ();
 sg13g2_decap_8 FILLER_12_1365 ();
 sg13g2_decap_8 FILLER_12_1372 ();
 sg13g2_decap_8 FILLER_12_1379 ();
 sg13g2_decap_8 FILLER_12_1386 ();
 sg13g2_decap_8 FILLER_12_1393 ();
 sg13g2_decap_8 FILLER_12_1400 ();
 sg13g2_decap_8 FILLER_12_1407 ();
 sg13g2_decap_8 FILLER_12_1414 ();
 sg13g2_decap_8 FILLER_12_1421 ();
 sg13g2_decap_8 FILLER_12_1428 ();
 sg13g2_decap_8 FILLER_12_1435 ();
 sg13g2_decap_8 FILLER_12_1442 ();
 sg13g2_decap_8 FILLER_12_1449 ();
 sg13g2_decap_8 FILLER_12_1456 ();
 sg13g2_decap_8 FILLER_12_1463 ();
 sg13g2_decap_8 FILLER_12_1470 ();
 sg13g2_decap_8 FILLER_12_1477 ();
 sg13g2_decap_8 FILLER_12_1484 ();
 sg13g2_decap_8 FILLER_12_1491 ();
 sg13g2_decap_8 FILLER_12_1498 ();
 sg13g2_decap_8 FILLER_12_1505 ();
 sg13g2_decap_8 FILLER_12_1512 ();
 sg13g2_decap_8 FILLER_12_1519 ();
 sg13g2_decap_8 FILLER_12_1526 ();
 sg13g2_decap_8 FILLER_12_1533 ();
 sg13g2_decap_8 FILLER_12_1540 ();
 sg13g2_decap_8 FILLER_12_1547 ();
 sg13g2_decap_8 FILLER_12_1554 ();
 sg13g2_decap_8 FILLER_12_1561 ();
 sg13g2_decap_8 FILLER_12_1568 ();
 sg13g2_decap_8 FILLER_12_1575 ();
 sg13g2_decap_8 FILLER_12_1582 ();
 sg13g2_decap_8 FILLER_12_1589 ();
 sg13g2_decap_8 FILLER_12_1596 ();
 sg13g2_decap_8 FILLER_12_1603 ();
 sg13g2_decap_8 FILLER_12_1610 ();
 sg13g2_decap_8 FILLER_12_1617 ();
 sg13g2_decap_8 FILLER_12_1624 ();
 sg13g2_decap_8 FILLER_12_1631 ();
 sg13g2_decap_8 FILLER_12_1638 ();
 sg13g2_decap_8 FILLER_12_1645 ();
 sg13g2_decap_8 FILLER_12_1652 ();
 sg13g2_decap_8 FILLER_12_1659 ();
 sg13g2_decap_8 FILLER_12_1666 ();
 sg13g2_decap_8 FILLER_12_1673 ();
 sg13g2_decap_8 FILLER_12_1680 ();
 sg13g2_decap_8 FILLER_12_1687 ();
 sg13g2_decap_8 FILLER_12_1694 ();
 sg13g2_decap_8 FILLER_12_1701 ();
 sg13g2_decap_8 FILLER_12_1708 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_decap_8 FILLER_12_1722 ();
 sg13g2_decap_8 FILLER_12_1729 ();
 sg13g2_decap_8 FILLER_12_1736 ();
 sg13g2_decap_8 FILLER_12_1743 ();
 sg13g2_decap_8 FILLER_12_1750 ();
 sg13g2_decap_8 FILLER_12_1757 ();
 sg13g2_decap_8 FILLER_12_1764 ();
 sg13g2_decap_8 FILLER_12_1771 ();
 sg13g2_decap_8 FILLER_12_1778 ();
 sg13g2_decap_8 FILLER_12_1785 ();
 sg13g2_decap_8 FILLER_12_1792 ();
 sg13g2_decap_8 FILLER_12_1799 ();
 sg13g2_decap_8 FILLER_12_1806 ();
 sg13g2_decap_8 FILLER_12_1813 ();
 sg13g2_decap_8 FILLER_12_1820 ();
 sg13g2_decap_8 FILLER_12_1827 ();
 sg13g2_decap_8 FILLER_12_1834 ();
 sg13g2_decap_8 FILLER_12_1841 ();
 sg13g2_decap_8 FILLER_12_1848 ();
 sg13g2_decap_8 FILLER_12_1855 ();
 sg13g2_decap_8 FILLER_12_1862 ();
 sg13g2_decap_8 FILLER_12_1869 ();
 sg13g2_decap_8 FILLER_12_1876 ();
 sg13g2_decap_8 FILLER_12_1883 ();
 sg13g2_decap_8 FILLER_12_1890 ();
 sg13g2_decap_8 FILLER_12_1897 ();
 sg13g2_decap_8 FILLER_12_1904 ();
 sg13g2_decap_8 FILLER_12_1911 ();
 sg13g2_decap_8 FILLER_12_1918 ();
 sg13g2_decap_8 FILLER_12_1925 ();
 sg13g2_decap_8 FILLER_12_1932 ();
 sg13g2_decap_8 FILLER_12_1939 ();
 sg13g2_decap_8 FILLER_12_1946 ();
 sg13g2_decap_8 FILLER_12_1953 ();
 sg13g2_decap_8 FILLER_12_1960 ();
 sg13g2_decap_8 FILLER_12_1967 ();
 sg13g2_decap_8 FILLER_12_1974 ();
 sg13g2_decap_8 FILLER_12_1981 ();
 sg13g2_decap_8 FILLER_12_1988 ();
 sg13g2_decap_8 FILLER_12_1995 ();
 sg13g2_decap_8 FILLER_12_2002 ();
 sg13g2_decap_8 FILLER_12_2009 ();
 sg13g2_decap_8 FILLER_12_2016 ();
 sg13g2_decap_8 FILLER_12_2023 ();
 sg13g2_decap_8 FILLER_12_2030 ();
 sg13g2_decap_8 FILLER_12_2037 ();
 sg13g2_decap_8 FILLER_12_2044 ();
 sg13g2_decap_8 FILLER_12_2051 ();
 sg13g2_fill_2 FILLER_12_2058 ();
 sg13g2_decap_8 FILLER_12_2081 ();
 sg13g2_decap_8 FILLER_12_2088 ();
 sg13g2_decap_8 FILLER_12_2095 ();
 sg13g2_decap_8 FILLER_12_2102 ();
 sg13g2_decap_8 FILLER_12_2109 ();
 sg13g2_decap_8 FILLER_12_2116 ();
 sg13g2_decap_8 FILLER_12_2123 ();
 sg13g2_decap_4 FILLER_12_2130 ();
 sg13g2_fill_1 FILLER_12_2134 ();
 sg13g2_decap_8 FILLER_12_2160 ();
 sg13g2_decap_4 FILLER_12_2167 ();
 sg13g2_decap_8 FILLER_12_2174 ();
 sg13g2_decap_8 FILLER_12_2181 ();
 sg13g2_decap_8 FILLER_12_2188 ();
 sg13g2_decap_8 FILLER_12_2195 ();
 sg13g2_decap_4 FILLER_12_2202 ();
 sg13g2_fill_2 FILLER_12_2206 ();
 sg13g2_decap_8 FILLER_12_2229 ();
 sg13g2_decap_8 FILLER_12_2236 ();
 sg13g2_decap_8 FILLER_12_2243 ();
 sg13g2_decap_8 FILLER_12_2250 ();
 sg13g2_decap_4 FILLER_12_2257 ();
 sg13g2_fill_1 FILLER_12_2261 ();
 sg13g2_decap_8 FILLER_12_2277 ();
 sg13g2_decap_8 FILLER_12_2284 ();
 sg13g2_decap_8 FILLER_12_2291 ();
 sg13g2_decap_8 FILLER_12_2298 ();
 sg13g2_decap_8 FILLER_12_2305 ();
 sg13g2_decap_8 FILLER_12_2312 ();
 sg13g2_decap_8 FILLER_12_2319 ();
 sg13g2_decap_8 FILLER_12_2326 ();
 sg13g2_decap_8 FILLER_12_2333 ();
 sg13g2_decap_8 FILLER_12_2340 ();
 sg13g2_decap_8 FILLER_12_2347 ();
 sg13g2_decap_8 FILLER_12_2359 ();
 sg13g2_decap_8 FILLER_12_2366 ();
 sg13g2_decap_8 FILLER_12_2373 ();
 sg13g2_decap_8 FILLER_12_2380 ();
 sg13g2_decap_8 FILLER_12_2387 ();
 sg13g2_decap_8 FILLER_12_2394 ();
 sg13g2_decap_8 FILLER_12_2401 ();
 sg13g2_fill_1 FILLER_12_2408 ();
 sg13g2_decap_8 FILLER_12_2434 ();
 sg13g2_decap_8 FILLER_12_2441 ();
 sg13g2_decap_8 FILLER_12_2448 ();
 sg13g2_decap_8 FILLER_12_2455 ();
 sg13g2_decap_8 FILLER_12_2462 ();
 sg13g2_decap_8 FILLER_12_2469 ();
 sg13g2_decap_8 FILLER_12_2476 ();
 sg13g2_decap_8 FILLER_12_2483 ();
 sg13g2_decap_8 FILLER_12_2490 ();
 sg13g2_decap_8 FILLER_12_2522 ();
 sg13g2_decap_8 FILLER_12_2529 ();
 sg13g2_decap_8 FILLER_12_2536 ();
 sg13g2_decap_8 FILLER_12_2543 ();
 sg13g2_fill_1 FILLER_12_2550 ();
 sg13g2_decap_8 FILLER_12_2564 ();
 sg13g2_decap_8 FILLER_12_2571 ();
 sg13g2_fill_2 FILLER_12_2578 ();
 sg13g2_decap_4 FILLER_12_2586 ();
 sg13g2_fill_2 FILLER_12_2590 ();
 sg13g2_decap_8 FILLER_12_2598 ();
 sg13g2_decap_8 FILLER_12_2605 ();
 sg13g2_decap_4 FILLER_12_2612 ();
 sg13g2_fill_1 FILLER_12_2616 ();
 sg13g2_decap_8 FILLER_12_2630 ();
 sg13g2_decap_8 FILLER_12_2637 ();
 sg13g2_decap_8 FILLER_12_2644 ();
 sg13g2_fill_1 FILLER_12_2651 ();
 sg13g2_fill_1 FILLER_12_2663 ();
 sg13g2_decap_8 FILLER_12_2667 ();
 sg13g2_fill_1 FILLER_12_2674 ();
 sg13g2_decap_8 FILLER_12_2688 ();
 sg13g2_decap_4 FILLER_12_2695 ();
 sg13g2_fill_1 FILLER_12_2699 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_fill_2 FILLER_13_560 ();
 sg13g2_fill_1 FILLER_13_562 ();
 sg13g2_decap_8 FILLER_13_584 ();
 sg13g2_decap_8 FILLER_13_591 ();
 sg13g2_decap_8 FILLER_13_598 ();
 sg13g2_decap_8 FILLER_13_605 ();
 sg13g2_decap_8 FILLER_13_633 ();
 sg13g2_decap_8 FILLER_13_640 ();
 sg13g2_decap_8 FILLER_13_647 ();
 sg13g2_fill_2 FILLER_13_654 ();
 sg13g2_decap_8 FILLER_13_677 ();
 sg13g2_decap_8 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_691 ();
 sg13g2_decap_4 FILLER_13_698 ();
 sg13g2_decap_8 FILLER_13_723 ();
 sg13g2_decap_8 FILLER_13_730 ();
 sg13g2_decap_8 FILLER_13_737 ();
 sg13g2_decap_8 FILLER_13_744 ();
 sg13g2_decap_8 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_758 ();
 sg13g2_fill_2 FILLER_13_765 ();
 sg13g2_decap_4 FILLER_13_792 ();
 sg13g2_decap_8 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_decap_8 FILLER_13_835 ();
 sg13g2_decap_8 FILLER_13_842 ();
 sg13g2_decap_8 FILLER_13_849 ();
 sg13g2_decap_8 FILLER_13_856 ();
 sg13g2_decap_8 FILLER_13_863 ();
 sg13g2_decap_8 FILLER_13_870 ();
 sg13g2_decap_8 FILLER_13_877 ();
 sg13g2_decap_8 FILLER_13_884 ();
 sg13g2_fill_2 FILLER_13_891 ();
 sg13g2_fill_1 FILLER_13_893 ();
 sg13g2_decap_8 FILLER_13_919 ();
 sg13g2_decap_8 FILLER_13_926 ();
 sg13g2_decap_8 FILLER_13_933 ();
 sg13g2_decap_8 FILLER_13_940 ();
 sg13g2_decap_8 FILLER_13_947 ();
 sg13g2_decap_8 FILLER_13_954 ();
 sg13g2_decap_8 FILLER_13_961 ();
 sg13g2_decap_8 FILLER_13_968 ();
 sg13g2_decap_8 FILLER_13_975 ();
 sg13g2_fill_2 FILLER_13_982 ();
 sg13g2_decap_8 FILLER_13_993 ();
 sg13g2_decap_8 FILLER_13_1000 ();
 sg13g2_decap_8 FILLER_13_1007 ();
 sg13g2_decap_8 FILLER_13_1014 ();
 sg13g2_decap_8 FILLER_13_1021 ();
 sg13g2_decap_8 FILLER_13_1028 ();
 sg13g2_decap_8 FILLER_13_1035 ();
 sg13g2_decap_8 FILLER_13_1042 ();
 sg13g2_decap_8 FILLER_13_1049 ();
 sg13g2_decap_8 FILLER_13_1056 ();
 sg13g2_decap_8 FILLER_13_1063 ();
 sg13g2_decap_8 FILLER_13_1070 ();
 sg13g2_decap_8 FILLER_13_1077 ();
 sg13g2_decap_8 FILLER_13_1084 ();
 sg13g2_decap_8 FILLER_13_1091 ();
 sg13g2_decap_8 FILLER_13_1098 ();
 sg13g2_decap_8 FILLER_13_1105 ();
 sg13g2_decap_8 FILLER_13_1112 ();
 sg13g2_decap_8 FILLER_13_1119 ();
 sg13g2_decap_8 FILLER_13_1126 ();
 sg13g2_decap_8 FILLER_13_1133 ();
 sg13g2_fill_2 FILLER_13_1140 ();
 sg13g2_fill_1 FILLER_13_1142 ();
 sg13g2_decap_8 FILLER_13_1168 ();
 sg13g2_decap_8 FILLER_13_1175 ();
 sg13g2_decap_8 FILLER_13_1182 ();
 sg13g2_decap_8 FILLER_13_1189 ();
 sg13g2_decap_8 FILLER_13_1196 ();
 sg13g2_decap_8 FILLER_13_1203 ();
 sg13g2_decap_8 FILLER_13_1210 ();
 sg13g2_decap_8 FILLER_13_1217 ();
 sg13g2_decap_8 FILLER_13_1224 ();
 sg13g2_decap_8 FILLER_13_1231 ();
 sg13g2_decap_8 FILLER_13_1238 ();
 sg13g2_decap_8 FILLER_13_1245 ();
 sg13g2_decap_8 FILLER_13_1252 ();
 sg13g2_decap_8 FILLER_13_1259 ();
 sg13g2_decap_8 FILLER_13_1266 ();
 sg13g2_decap_8 FILLER_13_1273 ();
 sg13g2_fill_2 FILLER_13_1280 ();
 sg13g2_fill_1 FILLER_13_1282 ();
 sg13g2_decap_8 FILLER_13_1308 ();
 sg13g2_decap_8 FILLER_13_1315 ();
 sg13g2_decap_8 FILLER_13_1322 ();
 sg13g2_fill_2 FILLER_13_1329 ();
 sg13g2_decap_8 FILLER_13_1336 ();
 sg13g2_decap_8 FILLER_13_1343 ();
 sg13g2_decap_8 FILLER_13_1350 ();
 sg13g2_decap_8 FILLER_13_1357 ();
 sg13g2_decap_8 FILLER_13_1364 ();
 sg13g2_decap_8 FILLER_13_1371 ();
 sg13g2_decap_8 FILLER_13_1378 ();
 sg13g2_decap_8 FILLER_13_1385 ();
 sg13g2_decap_8 FILLER_13_1392 ();
 sg13g2_decap_8 FILLER_13_1399 ();
 sg13g2_decap_8 FILLER_13_1406 ();
 sg13g2_decap_8 FILLER_13_1413 ();
 sg13g2_decap_8 FILLER_13_1420 ();
 sg13g2_decap_8 FILLER_13_1427 ();
 sg13g2_decap_8 FILLER_13_1434 ();
 sg13g2_decap_8 FILLER_13_1441 ();
 sg13g2_decap_8 FILLER_13_1448 ();
 sg13g2_decap_8 FILLER_13_1455 ();
 sg13g2_decap_8 FILLER_13_1462 ();
 sg13g2_fill_2 FILLER_13_1469 ();
 sg13g2_decap_8 FILLER_13_1474 ();
 sg13g2_decap_8 FILLER_13_1481 ();
 sg13g2_decap_8 FILLER_13_1488 ();
 sg13g2_decap_8 FILLER_13_1495 ();
 sg13g2_decap_8 FILLER_13_1502 ();
 sg13g2_decap_8 FILLER_13_1509 ();
 sg13g2_fill_1 FILLER_13_1516 ();
 sg13g2_decap_8 FILLER_13_1520 ();
 sg13g2_decap_8 FILLER_13_1527 ();
 sg13g2_decap_8 FILLER_13_1534 ();
 sg13g2_decap_8 FILLER_13_1541 ();
 sg13g2_decap_8 FILLER_13_1548 ();
 sg13g2_decap_8 FILLER_13_1555 ();
 sg13g2_decap_8 FILLER_13_1562 ();
 sg13g2_decap_8 FILLER_13_1569 ();
 sg13g2_decap_8 FILLER_13_1576 ();
 sg13g2_decap_8 FILLER_13_1583 ();
 sg13g2_decap_8 FILLER_13_1590 ();
 sg13g2_decap_8 FILLER_13_1600 ();
 sg13g2_decap_8 FILLER_13_1607 ();
 sg13g2_decap_8 FILLER_13_1614 ();
 sg13g2_decap_8 FILLER_13_1621 ();
 sg13g2_decap_8 FILLER_13_1628 ();
 sg13g2_decap_8 FILLER_13_1635 ();
 sg13g2_decap_8 FILLER_13_1642 ();
 sg13g2_decap_8 FILLER_13_1649 ();
 sg13g2_decap_8 FILLER_13_1656 ();
 sg13g2_decap_8 FILLER_13_1663 ();
 sg13g2_decap_8 FILLER_13_1670 ();
 sg13g2_decap_8 FILLER_13_1677 ();
 sg13g2_decap_8 FILLER_13_1684 ();
 sg13g2_decap_8 FILLER_13_1691 ();
 sg13g2_decap_8 FILLER_13_1698 ();
 sg13g2_decap_8 FILLER_13_1705 ();
 sg13g2_decap_8 FILLER_13_1712 ();
 sg13g2_decap_8 FILLER_13_1719 ();
 sg13g2_decap_8 FILLER_13_1726 ();
 sg13g2_decap_8 FILLER_13_1733 ();
 sg13g2_decap_8 FILLER_13_1740 ();
 sg13g2_decap_8 FILLER_13_1747 ();
 sg13g2_decap_8 FILLER_13_1754 ();
 sg13g2_decap_8 FILLER_13_1761 ();
 sg13g2_decap_8 FILLER_13_1768 ();
 sg13g2_decap_8 FILLER_13_1775 ();
 sg13g2_decap_8 FILLER_13_1782 ();
 sg13g2_decap_8 FILLER_13_1789 ();
 sg13g2_decap_8 FILLER_13_1796 ();
 sg13g2_decap_8 FILLER_13_1803 ();
 sg13g2_decap_8 FILLER_13_1810 ();
 sg13g2_decap_8 FILLER_13_1817 ();
 sg13g2_decap_8 FILLER_13_1824 ();
 sg13g2_decap_8 FILLER_13_1831 ();
 sg13g2_decap_8 FILLER_13_1838 ();
 sg13g2_decap_8 FILLER_13_1845 ();
 sg13g2_decap_8 FILLER_13_1852 ();
 sg13g2_decap_8 FILLER_13_1859 ();
 sg13g2_decap_8 FILLER_13_1866 ();
 sg13g2_decap_8 FILLER_13_1873 ();
 sg13g2_decap_8 FILLER_13_1880 ();
 sg13g2_decap_8 FILLER_13_1887 ();
 sg13g2_decap_8 FILLER_13_1894 ();
 sg13g2_decap_8 FILLER_13_1901 ();
 sg13g2_decap_4 FILLER_13_1908 ();
 sg13g2_decap_8 FILLER_13_1917 ();
 sg13g2_decap_8 FILLER_13_1924 ();
 sg13g2_decap_8 FILLER_13_1931 ();
 sg13g2_decap_8 FILLER_13_1938 ();
 sg13g2_decap_8 FILLER_13_1945 ();
 sg13g2_decap_8 FILLER_13_1952 ();
 sg13g2_decap_8 FILLER_13_1959 ();
 sg13g2_decap_8 FILLER_13_1966 ();
 sg13g2_decap_8 FILLER_13_1973 ();
 sg13g2_decap_8 FILLER_13_1980 ();
 sg13g2_decap_8 FILLER_13_1987 ();
 sg13g2_decap_8 FILLER_13_1994 ();
 sg13g2_decap_8 FILLER_13_2001 ();
 sg13g2_decap_8 FILLER_13_2008 ();
 sg13g2_decap_8 FILLER_13_2015 ();
 sg13g2_decap_8 FILLER_13_2022 ();
 sg13g2_decap_8 FILLER_13_2029 ();
 sg13g2_decap_8 FILLER_13_2036 ();
 sg13g2_decap_8 FILLER_13_2043 ();
 sg13g2_decap_4 FILLER_13_2050 ();
 sg13g2_decap_8 FILLER_13_2079 ();
 sg13g2_decap_8 FILLER_13_2086 ();
 sg13g2_decap_8 FILLER_13_2093 ();
 sg13g2_decap_8 FILLER_13_2100 ();
 sg13g2_fill_2 FILLER_13_2107 ();
 sg13g2_decap_8 FILLER_13_2112 ();
 sg13g2_decap_8 FILLER_13_2119 ();
 sg13g2_decap_8 FILLER_13_2126 ();
 sg13g2_decap_8 FILLER_13_2133 ();
 sg13g2_decap_8 FILLER_13_2140 ();
 sg13g2_decap_8 FILLER_13_2147 ();
 sg13g2_decap_8 FILLER_13_2154 ();
 sg13g2_decap_8 FILLER_13_2161 ();
 sg13g2_decap_8 FILLER_13_2168 ();
 sg13g2_decap_8 FILLER_13_2175 ();
 sg13g2_decap_8 FILLER_13_2182 ();
 sg13g2_decap_8 FILLER_13_2189 ();
 sg13g2_decap_8 FILLER_13_2196 ();
 sg13g2_fill_2 FILLER_13_2203 ();
 sg13g2_decap_8 FILLER_13_2230 ();
 sg13g2_decap_8 FILLER_13_2237 ();
 sg13g2_decap_8 FILLER_13_2244 ();
 sg13g2_decap_8 FILLER_13_2251 ();
 sg13g2_decap_8 FILLER_13_2258 ();
 sg13g2_decap_8 FILLER_13_2265 ();
 sg13g2_decap_8 FILLER_13_2272 ();
 sg13g2_decap_8 FILLER_13_2279 ();
 sg13g2_decap_8 FILLER_13_2286 ();
 sg13g2_decap_8 FILLER_13_2293 ();
 sg13g2_decap_8 FILLER_13_2300 ();
 sg13g2_decap_8 FILLER_13_2307 ();
 sg13g2_decap_8 FILLER_13_2314 ();
 sg13g2_decap_4 FILLER_13_2321 ();
 sg13g2_fill_1 FILLER_13_2325 ();
 sg13g2_decap_8 FILLER_13_2341 ();
 sg13g2_decap_8 FILLER_13_2348 ();
 sg13g2_decap_8 FILLER_13_2355 ();
 sg13g2_decap_8 FILLER_13_2362 ();
 sg13g2_decap_8 FILLER_13_2369 ();
 sg13g2_decap_8 FILLER_13_2376 ();
 sg13g2_decap_8 FILLER_13_2383 ();
 sg13g2_decap_8 FILLER_13_2390 ();
 sg13g2_decap_8 FILLER_13_2397 ();
 sg13g2_decap_8 FILLER_13_2404 ();
 sg13g2_decap_8 FILLER_13_2411 ();
 sg13g2_fill_2 FILLER_13_2418 ();
 sg13g2_decap_8 FILLER_13_2425 ();
 sg13g2_decap_8 FILLER_13_2432 ();
 sg13g2_decap_8 FILLER_13_2439 ();
 sg13g2_decap_8 FILLER_13_2446 ();
 sg13g2_decap_8 FILLER_13_2453 ();
 sg13g2_decap_8 FILLER_13_2460 ();
 sg13g2_decap_4 FILLER_13_2467 ();
 sg13g2_fill_1 FILLER_13_2471 ();
 sg13g2_decap_8 FILLER_13_2488 ();
 sg13g2_decap_8 FILLER_13_2495 ();
 sg13g2_decap_8 FILLER_13_2502 ();
 sg13g2_decap_8 FILLER_13_2509 ();
 sg13g2_decap_8 FILLER_13_2516 ();
 sg13g2_decap_8 FILLER_13_2523 ();
 sg13g2_decap_8 FILLER_13_2530 ();
 sg13g2_decap_8 FILLER_13_2537 ();
 sg13g2_decap_8 FILLER_13_2544 ();
 sg13g2_decap_8 FILLER_13_2551 ();
 sg13g2_decap_8 FILLER_13_2558 ();
 sg13g2_decap_8 FILLER_13_2565 ();
 sg13g2_fill_2 FILLER_13_2572 ();
 sg13g2_fill_1 FILLER_13_2574 ();
 sg13g2_decap_8 FILLER_13_2601 ();
 sg13g2_decap_8 FILLER_13_2608 ();
 sg13g2_decap_8 FILLER_13_2615 ();
 sg13g2_decap_8 FILLER_13_2622 ();
 sg13g2_decap_8 FILLER_13_2629 ();
 sg13g2_decap_8 FILLER_13_2636 ();
 sg13g2_decap_8 FILLER_13_2643 ();
 sg13g2_fill_2 FILLER_13_2650 ();
 sg13g2_decap_8 FILLER_13_2662 ();
 sg13g2_fill_2 FILLER_13_2669 ();
 sg13g2_decap_4 FILLER_13_2676 ();
 sg13g2_fill_1 FILLER_13_2680 ();
 sg13g2_decap_8 FILLER_13_2689 ();
 sg13g2_decap_4 FILLER_13_2696 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_4 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_430 ();
 sg13g2_decap_8 FILLER_14_437 ();
 sg13g2_decap_8 FILLER_14_444 ();
 sg13g2_decap_8 FILLER_14_451 ();
 sg13g2_decap_8 FILLER_14_458 ();
 sg13g2_decap_8 FILLER_14_465 ();
 sg13g2_decap_8 FILLER_14_472 ();
 sg13g2_decap_8 FILLER_14_479 ();
 sg13g2_decap_8 FILLER_14_486 ();
 sg13g2_decap_8 FILLER_14_493 ();
 sg13g2_decap_8 FILLER_14_500 ();
 sg13g2_decap_8 FILLER_14_507 ();
 sg13g2_decap_8 FILLER_14_514 ();
 sg13g2_decap_8 FILLER_14_521 ();
 sg13g2_decap_8 FILLER_14_528 ();
 sg13g2_decap_8 FILLER_14_535 ();
 sg13g2_decap_8 FILLER_14_542 ();
 sg13g2_decap_8 FILLER_14_549 ();
 sg13g2_decap_8 FILLER_14_556 ();
 sg13g2_decap_8 FILLER_14_563 ();
 sg13g2_decap_8 FILLER_14_570 ();
 sg13g2_decap_8 FILLER_14_577 ();
 sg13g2_decap_8 FILLER_14_584 ();
 sg13g2_decap_8 FILLER_14_591 ();
 sg13g2_decap_8 FILLER_14_598 ();
 sg13g2_decap_8 FILLER_14_605 ();
 sg13g2_decap_8 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_619 ();
 sg13g2_decap_8 FILLER_14_626 ();
 sg13g2_decap_8 FILLER_14_633 ();
 sg13g2_decap_8 FILLER_14_640 ();
 sg13g2_decap_4 FILLER_14_647 ();
 sg13g2_fill_2 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_656 ();
 sg13g2_decap_8 FILLER_14_663 ();
 sg13g2_decap_8 FILLER_14_670 ();
 sg13g2_decap_8 FILLER_14_677 ();
 sg13g2_decap_8 FILLER_14_684 ();
 sg13g2_decap_8 FILLER_14_691 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_decap_8 FILLER_14_705 ();
 sg13g2_decap_8 FILLER_14_712 ();
 sg13g2_decap_8 FILLER_14_719 ();
 sg13g2_decap_8 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_733 ();
 sg13g2_decap_8 FILLER_14_740 ();
 sg13g2_decap_8 FILLER_14_747 ();
 sg13g2_decap_8 FILLER_14_754 ();
 sg13g2_decap_8 FILLER_14_761 ();
 sg13g2_decap_8 FILLER_14_768 ();
 sg13g2_decap_8 FILLER_14_775 ();
 sg13g2_decap_8 FILLER_14_782 ();
 sg13g2_decap_8 FILLER_14_789 ();
 sg13g2_decap_8 FILLER_14_796 ();
 sg13g2_decap_8 FILLER_14_803 ();
 sg13g2_decap_8 FILLER_14_810 ();
 sg13g2_decap_8 FILLER_14_817 ();
 sg13g2_decap_8 FILLER_14_824 ();
 sg13g2_decap_8 FILLER_14_831 ();
 sg13g2_decap_8 FILLER_14_838 ();
 sg13g2_decap_8 FILLER_14_845 ();
 sg13g2_decap_8 FILLER_14_852 ();
 sg13g2_decap_8 FILLER_14_859 ();
 sg13g2_fill_2 FILLER_14_866 ();
 sg13g2_fill_1 FILLER_14_868 ();
 sg13g2_decap_8 FILLER_14_882 ();
 sg13g2_decap_8 FILLER_14_889 ();
 sg13g2_decap_8 FILLER_14_896 ();
 sg13g2_decap_8 FILLER_14_903 ();
 sg13g2_decap_8 FILLER_14_910 ();
 sg13g2_decap_8 FILLER_14_917 ();
 sg13g2_decap_4 FILLER_14_924 ();
 sg13g2_fill_2 FILLER_14_928 ();
 sg13g2_decap_8 FILLER_14_955 ();
 sg13g2_decap_8 FILLER_14_962 ();
 sg13g2_decap_4 FILLER_14_969 ();
 sg13g2_decap_8 FILLER_14_983 ();
 sg13g2_fill_1 FILLER_14_990 ();
 sg13g2_decap_8 FILLER_14_996 ();
 sg13g2_decap_8 FILLER_14_1003 ();
 sg13g2_decap_8 FILLER_14_1010 ();
 sg13g2_decap_8 FILLER_14_1017 ();
 sg13g2_decap_8 FILLER_14_1024 ();
 sg13g2_fill_1 FILLER_14_1031 ();
 sg13g2_decap_8 FILLER_14_1053 ();
 sg13g2_decap_8 FILLER_14_1060 ();
 sg13g2_decap_8 FILLER_14_1067 ();
 sg13g2_decap_4 FILLER_14_1074 ();
 sg13g2_fill_2 FILLER_14_1078 ();
 sg13g2_decap_8 FILLER_14_1101 ();
 sg13g2_decap_8 FILLER_14_1108 ();
 sg13g2_decap_8 FILLER_14_1115 ();
 sg13g2_decap_8 FILLER_14_1122 ();
 sg13g2_decap_8 FILLER_14_1129 ();
 sg13g2_decap_8 FILLER_14_1136 ();
 sg13g2_decap_8 FILLER_14_1143 ();
 sg13g2_fill_2 FILLER_14_1150 ();
 sg13g2_fill_1 FILLER_14_1152 ();
 sg13g2_decap_8 FILLER_14_1174 ();
 sg13g2_decap_8 FILLER_14_1181 ();
 sg13g2_decap_8 FILLER_14_1188 ();
 sg13g2_decap_8 FILLER_14_1195 ();
 sg13g2_decap_8 FILLER_14_1202 ();
 sg13g2_decap_8 FILLER_14_1209 ();
 sg13g2_decap_8 FILLER_14_1216 ();
 sg13g2_decap_8 FILLER_14_1223 ();
 sg13g2_decap_8 FILLER_14_1230 ();
 sg13g2_decap_8 FILLER_14_1237 ();
 sg13g2_decap_8 FILLER_14_1244 ();
 sg13g2_decap_8 FILLER_14_1251 ();
 sg13g2_decap_8 FILLER_14_1258 ();
 sg13g2_decap_8 FILLER_14_1265 ();
 sg13g2_decap_8 FILLER_14_1272 ();
 sg13g2_decap_8 FILLER_14_1279 ();
 sg13g2_decap_8 FILLER_14_1286 ();
 sg13g2_decap_8 FILLER_14_1293 ();
 sg13g2_decap_8 FILLER_14_1300 ();
 sg13g2_decap_8 FILLER_14_1307 ();
 sg13g2_decap_8 FILLER_14_1314 ();
 sg13g2_decap_8 FILLER_14_1321 ();
 sg13g2_decap_8 FILLER_14_1341 ();
 sg13g2_decap_8 FILLER_14_1348 ();
 sg13g2_decap_8 FILLER_14_1355 ();
 sg13g2_decap_8 FILLER_14_1362 ();
 sg13g2_decap_8 FILLER_14_1369 ();
 sg13g2_decap_8 FILLER_14_1376 ();
 sg13g2_decap_8 FILLER_14_1383 ();
 sg13g2_decap_8 FILLER_14_1390 ();
 sg13g2_decap_8 FILLER_14_1397 ();
 sg13g2_decap_8 FILLER_14_1404 ();
 sg13g2_decap_8 FILLER_14_1411 ();
 sg13g2_decap_8 FILLER_14_1418 ();
 sg13g2_decap_8 FILLER_14_1425 ();
 sg13g2_decap_8 FILLER_14_1432 ();
 sg13g2_decap_8 FILLER_14_1439 ();
 sg13g2_decap_8 FILLER_14_1446 ();
 sg13g2_decap_8 FILLER_14_1453 ();
 sg13g2_decap_8 FILLER_14_1460 ();
 sg13g2_decap_8 FILLER_14_1467 ();
 sg13g2_decap_8 FILLER_14_1474 ();
 sg13g2_decap_8 FILLER_14_1481 ();
 sg13g2_decap_8 FILLER_14_1488 ();
 sg13g2_decap_8 FILLER_14_1495 ();
 sg13g2_decap_8 FILLER_14_1502 ();
 sg13g2_decap_8 FILLER_14_1509 ();
 sg13g2_decap_8 FILLER_14_1516 ();
 sg13g2_decap_8 FILLER_14_1523 ();
 sg13g2_decap_8 FILLER_14_1530 ();
 sg13g2_decap_8 FILLER_14_1537 ();
 sg13g2_decap_8 FILLER_14_1544 ();
 sg13g2_decap_8 FILLER_14_1551 ();
 sg13g2_decap_8 FILLER_14_1558 ();
 sg13g2_decap_8 FILLER_14_1565 ();
 sg13g2_decap_8 FILLER_14_1572 ();
 sg13g2_decap_8 FILLER_14_1579 ();
 sg13g2_decap_8 FILLER_14_1586 ();
 sg13g2_decap_8 FILLER_14_1593 ();
 sg13g2_decap_8 FILLER_14_1600 ();
 sg13g2_decap_8 FILLER_14_1607 ();
 sg13g2_decap_8 FILLER_14_1614 ();
 sg13g2_decap_8 FILLER_14_1621 ();
 sg13g2_decap_8 FILLER_14_1628 ();
 sg13g2_decap_8 FILLER_14_1635 ();
 sg13g2_decap_8 FILLER_14_1642 ();
 sg13g2_decap_8 FILLER_14_1649 ();
 sg13g2_decap_8 FILLER_14_1656 ();
 sg13g2_decap_8 FILLER_14_1663 ();
 sg13g2_decap_8 FILLER_14_1670 ();
 sg13g2_decap_8 FILLER_14_1677 ();
 sg13g2_decap_8 FILLER_14_1684 ();
 sg13g2_decap_8 FILLER_14_1691 ();
 sg13g2_decap_8 FILLER_14_1698 ();
 sg13g2_decap_8 FILLER_14_1705 ();
 sg13g2_decap_8 FILLER_14_1712 ();
 sg13g2_decap_8 FILLER_14_1719 ();
 sg13g2_decap_8 FILLER_14_1726 ();
 sg13g2_decap_8 FILLER_14_1733 ();
 sg13g2_decap_4 FILLER_14_1740 ();
 sg13g2_decap_8 FILLER_14_1767 ();
 sg13g2_decap_8 FILLER_14_1774 ();
 sg13g2_decap_8 FILLER_14_1781 ();
 sg13g2_decap_4 FILLER_14_1788 ();
 sg13g2_fill_2 FILLER_14_1792 ();
 sg13g2_fill_1 FILLER_14_1799 ();
 sg13g2_decap_8 FILLER_14_1813 ();
 sg13g2_decap_8 FILLER_14_1820 ();
 sg13g2_decap_8 FILLER_14_1827 ();
 sg13g2_decap_8 FILLER_14_1834 ();
 sg13g2_decap_8 FILLER_14_1841 ();
 sg13g2_decap_8 FILLER_14_1848 ();
 sg13g2_decap_8 FILLER_14_1855 ();
 sg13g2_decap_8 FILLER_14_1862 ();
 sg13g2_decap_8 FILLER_14_1869 ();
 sg13g2_decap_8 FILLER_14_1876 ();
 sg13g2_decap_8 FILLER_14_1883 ();
 sg13g2_decap_8 FILLER_14_1890 ();
 sg13g2_decap_8 FILLER_14_1897 ();
 sg13g2_decap_8 FILLER_14_1904 ();
 sg13g2_decap_8 FILLER_14_1911 ();
 sg13g2_decap_8 FILLER_14_1918 ();
 sg13g2_decap_8 FILLER_14_1925 ();
 sg13g2_decap_4 FILLER_14_1932 ();
 sg13g2_decap_8 FILLER_14_1957 ();
 sg13g2_decap_8 FILLER_14_1964 ();
 sg13g2_decap_8 FILLER_14_1971 ();
 sg13g2_decap_8 FILLER_14_1978 ();
 sg13g2_decap_4 FILLER_14_1985 ();
 sg13g2_fill_1 FILLER_14_1989 ();
 sg13g2_decap_8 FILLER_14_2011 ();
 sg13g2_decap_8 FILLER_14_2018 ();
 sg13g2_decap_8 FILLER_14_2025 ();
 sg13g2_decap_8 FILLER_14_2032 ();
 sg13g2_decap_8 FILLER_14_2039 ();
 sg13g2_decap_8 FILLER_14_2046 ();
 sg13g2_decap_8 FILLER_14_2053 ();
 sg13g2_decap_8 FILLER_14_2060 ();
 sg13g2_decap_8 FILLER_14_2067 ();
 sg13g2_decap_8 FILLER_14_2074 ();
 sg13g2_decap_8 FILLER_14_2081 ();
 sg13g2_decap_8 FILLER_14_2088 ();
 sg13g2_decap_8 FILLER_14_2095 ();
 sg13g2_decap_8 FILLER_14_2102 ();
 sg13g2_decap_8 FILLER_14_2109 ();
 sg13g2_decap_8 FILLER_14_2116 ();
 sg13g2_decap_8 FILLER_14_2123 ();
 sg13g2_decap_8 FILLER_14_2130 ();
 sg13g2_decap_8 FILLER_14_2137 ();
 sg13g2_decap_8 FILLER_14_2144 ();
 sg13g2_decap_8 FILLER_14_2151 ();
 sg13g2_decap_8 FILLER_14_2158 ();
 sg13g2_decap_8 FILLER_14_2165 ();
 sg13g2_decap_8 FILLER_14_2172 ();
 sg13g2_decap_8 FILLER_14_2179 ();
 sg13g2_decap_8 FILLER_14_2186 ();
 sg13g2_decap_8 FILLER_14_2193 ();
 sg13g2_decap_8 FILLER_14_2200 ();
 sg13g2_decap_8 FILLER_14_2207 ();
 sg13g2_decap_8 FILLER_14_2214 ();
 sg13g2_decap_8 FILLER_14_2221 ();
 sg13g2_decap_8 FILLER_14_2228 ();
 sg13g2_decap_8 FILLER_14_2245 ();
 sg13g2_decap_4 FILLER_14_2252 ();
 sg13g2_fill_1 FILLER_14_2256 ();
 sg13g2_decap_8 FILLER_14_2262 ();
 sg13g2_decap_8 FILLER_14_2269 ();
 sg13g2_decap_8 FILLER_14_2276 ();
 sg13g2_decap_8 FILLER_14_2283 ();
 sg13g2_decap_4 FILLER_14_2290 ();
 sg13g2_decap_8 FILLER_14_2309 ();
 sg13g2_decap_8 FILLER_14_2316 ();
 sg13g2_fill_2 FILLER_14_2323 ();
 sg13g2_fill_1 FILLER_14_2325 ();
 sg13g2_decap_8 FILLER_14_2341 ();
 sg13g2_decap_8 FILLER_14_2348 ();
 sg13g2_decap_8 FILLER_14_2355 ();
 sg13g2_decap_8 FILLER_14_2362 ();
 sg13g2_decap_8 FILLER_14_2369 ();
 sg13g2_decap_8 FILLER_14_2376 ();
 sg13g2_decap_4 FILLER_14_2383 ();
 sg13g2_decap_8 FILLER_14_2397 ();
 sg13g2_decap_8 FILLER_14_2404 ();
 sg13g2_fill_2 FILLER_14_2411 ();
 sg13g2_decap_8 FILLER_14_2416 ();
 sg13g2_decap_8 FILLER_14_2423 ();
 sg13g2_decap_8 FILLER_14_2430 ();
 sg13g2_decap_8 FILLER_14_2440 ();
 sg13g2_decap_8 FILLER_14_2447 ();
 sg13g2_fill_2 FILLER_14_2454 ();
 sg13g2_decap_8 FILLER_14_2459 ();
 sg13g2_decap_8 FILLER_14_2466 ();
 sg13g2_decap_8 FILLER_14_2473 ();
 sg13g2_fill_2 FILLER_14_2480 ();
 sg13g2_fill_1 FILLER_14_2482 ();
 sg13g2_decap_8 FILLER_14_2488 ();
 sg13g2_decap_8 FILLER_14_2495 ();
 sg13g2_decap_8 FILLER_14_2502 ();
 sg13g2_decap_4 FILLER_14_2509 ();
 sg13g2_fill_1 FILLER_14_2513 ();
 sg13g2_decap_8 FILLER_14_2519 ();
 sg13g2_decap_8 FILLER_14_2526 ();
 sg13g2_decap_4 FILLER_14_2533 ();
 sg13g2_fill_2 FILLER_14_2537 ();
 sg13g2_decap_8 FILLER_14_2555 ();
 sg13g2_decap_8 FILLER_14_2562 ();
 sg13g2_decap_8 FILLER_14_2569 ();
 sg13g2_decap_8 FILLER_14_2576 ();
 sg13g2_decap_8 FILLER_14_2583 ();
 sg13g2_decap_8 FILLER_14_2590 ();
 sg13g2_decap_8 FILLER_14_2597 ();
 sg13g2_decap_8 FILLER_14_2604 ();
 sg13g2_decap_8 FILLER_14_2611 ();
 sg13g2_decap_4 FILLER_14_2618 ();
 sg13g2_decap_8 FILLER_14_2635 ();
 sg13g2_decap_8 FILLER_14_2642 ();
 sg13g2_decap_8 FILLER_14_2649 ();
 sg13g2_decap_8 FILLER_14_2656 ();
 sg13g2_decap_4 FILLER_14_2663 ();
 sg13g2_fill_2 FILLER_14_2672 ();
 sg13g2_decap_4 FILLER_14_2696 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_fill_2 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_decap_8 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_15_414 ();
 sg13g2_decap_8 FILLER_15_421 ();
 sg13g2_decap_8 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_15_435 ();
 sg13g2_decap_8 FILLER_15_442 ();
 sg13g2_decap_8 FILLER_15_449 ();
 sg13g2_decap_8 FILLER_15_456 ();
 sg13g2_decap_8 FILLER_15_463 ();
 sg13g2_decap_8 FILLER_15_470 ();
 sg13g2_decap_8 FILLER_15_477 ();
 sg13g2_decap_8 FILLER_15_484 ();
 sg13g2_decap_8 FILLER_15_491 ();
 sg13g2_decap_8 FILLER_15_498 ();
 sg13g2_decap_8 FILLER_15_505 ();
 sg13g2_decap_8 FILLER_15_512 ();
 sg13g2_decap_8 FILLER_15_519 ();
 sg13g2_decap_8 FILLER_15_526 ();
 sg13g2_decap_8 FILLER_15_533 ();
 sg13g2_decap_8 FILLER_15_540 ();
 sg13g2_decap_8 FILLER_15_547 ();
 sg13g2_decap_8 FILLER_15_554 ();
 sg13g2_decap_8 FILLER_15_561 ();
 sg13g2_decap_8 FILLER_15_568 ();
 sg13g2_decap_8 FILLER_15_575 ();
 sg13g2_decap_8 FILLER_15_582 ();
 sg13g2_decap_8 FILLER_15_589 ();
 sg13g2_decap_8 FILLER_15_596 ();
 sg13g2_decap_4 FILLER_15_603 ();
 sg13g2_fill_2 FILLER_15_607 ();
 sg13g2_decap_8 FILLER_15_612 ();
 sg13g2_decap_8 FILLER_15_619 ();
 sg13g2_decap_8 FILLER_15_626 ();
 sg13g2_decap_8 FILLER_15_633 ();
 sg13g2_decap_8 FILLER_15_640 ();
 sg13g2_decap_8 FILLER_15_647 ();
 sg13g2_decap_8 FILLER_15_654 ();
 sg13g2_decap_8 FILLER_15_661 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_decap_8 FILLER_15_675 ();
 sg13g2_decap_8 FILLER_15_682 ();
 sg13g2_decap_8 FILLER_15_689 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_710 ();
 sg13g2_decap_8 FILLER_15_717 ();
 sg13g2_decap_8 FILLER_15_730 ();
 sg13g2_decap_8 FILLER_15_737 ();
 sg13g2_decap_8 FILLER_15_744 ();
 sg13g2_decap_8 FILLER_15_751 ();
 sg13g2_decap_8 FILLER_15_758 ();
 sg13g2_decap_8 FILLER_15_765 ();
 sg13g2_decap_8 FILLER_15_772 ();
 sg13g2_decap_8 FILLER_15_779 ();
 sg13g2_decap_8 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_793 ();
 sg13g2_decap_8 FILLER_15_800 ();
 sg13g2_decap_8 FILLER_15_807 ();
 sg13g2_decap_8 FILLER_15_814 ();
 sg13g2_decap_8 FILLER_15_821 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_decap_8 FILLER_15_835 ();
 sg13g2_decap_8 FILLER_15_842 ();
 sg13g2_decap_8 FILLER_15_849 ();
 sg13g2_decap_8 FILLER_15_856 ();
 sg13g2_decap_8 FILLER_15_863 ();
 sg13g2_decap_8 FILLER_15_870 ();
 sg13g2_decap_8 FILLER_15_877 ();
 sg13g2_decap_8 FILLER_15_884 ();
 sg13g2_decap_8 FILLER_15_891 ();
 sg13g2_decap_8 FILLER_15_898 ();
 sg13g2_decap_8 FILLER_15_905 ();
 sg13g2_decap_8 FILLER_15_912 ();
 sg13g2_decap_8 FILLER_15_919 ();
 sg13g2_decap_8 FILLER_15_926 ();
 sg13g2_decap_8 FILLER_15_933 ();
 sg13g2_decap_8 FILLER_15_940 ();
 sg13g2_decap_8 FILLER_15_947 ();
 sg13g2_decap_8 FILLER_15_954 ();
 sg13g2_decap_8 FILLER_15_961 ();
 sg13g2_decap_8 FILLER_15_968 ();
 sg13g2_decap_8 FILLER_15_975 ();
 sg13g2_decap_8 FILLER_15_982 ();
 sg13g2_decap_8 FILLER_15_989 ();
 sg13g2_decap_8 FILLER_15_996 ();
 sg13g2_decap_8 FILLER_15_1003 ();
 sg13g2_decap_8 FILLER_15_1010 ();
 sg13g2_decap_8 FILLER_15_1017 ();
 sg13g2_decap_4 FILLER_15_1024 ();
 sg13g2_fill_1 FILLER_15_1028 ();
 sg13g2_decap_8 FILLER_15_1054 ();
 sg13g2_decap_8 FILLER_15_1061 ();
 sg13g2_decap_8 FILLER_15_1068 ();
 sg13g2_decap_8 FILLER_15_1100 ();
 sg13g2_decap_8 FILLER_15_1107 ();
 sg13g2_decap_8 FILLER_15_1114 ();
 sg13g2_fill_1 FILLER_15_1121 ();
 sg13g2_decap_8 FILLER_15_1125 ();
 sg13g2_decap_8 FILLER_15_1132 ();
 sg13g2_decap_8 FILLER_15_1139 ();
 sg13g2_decap_8 FILLER_15_1146 ();
 sg13g2_decap_8 FILLER_15_1153 ();
 sg13g2_decap_8 FILLER_15_1160 ();
 sg13g2_decap_8 FILLER_15_1167 ();
 sg13g2_decap_8 FILLER_15_1174 ();
 sg13g2_decap_8 FILLER_15_1181 ();
 sg13g2_decap_8 FILLER_15_1188 ();
 sg13g2_decap_4 FILLER_15_1198 ();
 sg13g2_fill_2 FILLER_15_1202 ();
 sg13g2_decap_8 FILLER_15_1207 ();
 sg13g2_decap_8 FILLER_15_1214 ();
 sg13g2_decap_8 FILLER_15_1221 ();
 sg13g2_fill_2 FILLER_15_1228 ();
 sg13g2_decap_8 FILLER_15_1233 ();
 sg13g2_decap_8 FILLER_15_1240 ();
 sg13g2_decap_4 FILLER_15_1247 ();
 sg13g2_decap_8 FILLER_15_1254 ();
 sg13g2_decap_8 FILLER_15_1261 ();
 sg13g2_decap_8 FILLER_15_1268 ();
 sg13g2_decap_8 FILLER_15_1275 ();
 sg13g2_decap_8 FILLER_15_1285 ();
 sg13g2_decap_8 FILLER_15_1292 ();
 sg13g2_decap_8 FILLER_15_1299 ();
 sg13g2_decap_8 FILLER_15_1306 ();
 sg13g2_decap_8 FILLER_15_1313 ();
 sg13g2_decap_8 FILLER_15_1320 ();
 sg13g2_decap_8 FILLER_15_1327 ();
 sg13g2_decap_8 FILLER_15_1334 ();
 sg13g2_decap_8 FILLER_15_1341 ();
 sg13g2_decap_8 FILLER_15_1348 ();
 sg13g2_decap_8 FILLER_15_1355 ();
 sg13g2_decap_8 FILLER_15_1362 ();
 sg13g2_decap_8 FILLER_15_1369 ();
 sg13g2_decap_8 FILLER_15_1376 ();
 sg13g2_decap_8 FILLER_15_1383 ();
 sg13g2_decap_8 FILLER_15_1390 ();
 sg13g2_decap_8 FILLER_15_1397 ();
 sg13g2_decap_8 FILLER_15_1404 ();
 sg13g2_decap_8 FILLER_15_1411 ();
 sg13g2_decap_8 FILLER_15_1418 ();
 sg13g2_decap_8 FILLER_15_1425 ();
 sg13g2_decap_8 FILLER_15_1432 ();
 sg13g2_decap_8 FILLER_15_1439 ();
 sg13g2_decap_8 FILLER_15_1446 ();
 sg13g2_decap_8 FILLER_15_1453 ();
 sg13g2_decap_8 FILLER_15_1460 ();
 sg13g2_decap_8 FILLER_15_1467 ();
 sg13g2_decap_8 FILLER_15_1474 ();
 sg13g2_decap_8 FILLER_15_1481 ();
 sg13g2_decap_8 FILLER_15_1488 ();
 sg13g2_decap_8 FILLER_15_1495 ();
 sg13g2_decap_8 FILLER_15_1502 ();
 sg13g2_decap_8 FILLER_15_1509 ();
 sg13g2_decap_8 FILLER_15_1516 ();
 sg13g2_decap_8 FILLER_15_1523 ();
 sg13g2_decap_8 FILLER_15_1530 ();
 sg13g2_decap_8 FILLER_15_1537 ();
 sg13g2_decap_8 FILLER_15_1544 ();
 sg13g2_decap_8 FILLER_15_1551 ();
 sg13g2_decap_8 FILLER_15_1558 ();
 sg13g2_decap_8 FILLER_15_1565 ();
 sg13g2_decap_8 FILLER_15_1572 ();
 sg13g2_decap_8 FILLER_15_1579 ();
 sg13g2_decap_8 FILLER_15_1586 ();
 sg13g2_decap_8 FILLER_15_1593 ();
 sg13g2_decap_8 FILLER_15_1600 ();
 sg13g2_decap_8 FILLER_15_1607 ();
 sg13g2_decap_8 FILLER_15_1614 ();
 sg13g2_decap_8 FILLER_15_1621 ();
 sg13g2_decap_8 FILLER_15_1628 ();
 sg13g2_decap_8 FILLER_15_1635 ();
 sg13g2_decap_8 FILLER_15_1642 ();
 sg13g2_decap_8 FILLER_15_1649 ();
 sg13g2_decap_8 FILLER_15_1656 ();
 sg13g2_decap_8 FILLER_15_1663 ();
 sg13g2_decap_8 FILLER_15_1670 ();
 sg13g2_decap_8 FILLER_15_1677 ();
 sg13g2_decap_8 FILLER_15_1684 ();
 sg13g2_decap_8 FILLER_15_1691 ();
 sg13g2_decap_8 FILLER_15_1698 ();
 sg13g2_decap_8 FILLER_15_1705 ();
 sg13g2_decap_8 FILLER_15_1712 ();
 sg13g2_decap_8 FILLER_15_1719 ();
 sg13g2_decap_8 FILLER_15_1726 ();
 sg13g2_decap_8 FILLER_15_1733 ();
 sg13g2_decap_8 FILLER_15_1740 ();
 sg13g2_decap_8 FILLER_15_1747 ();
 sg13g2_decap_8 FILLER_15_1754 ();
 sg13g2_decap_8 FILLER_15_1761 ();
 sg13g2_decap_8 FILLER_15_1768 ();
 sg13g2_decap_8 FILLER_15_1775 ();
 sg13g2_decap_8 FILLER_15_1782 ();
 sg13g2_decap_8 FILLER_15_1789 ();
 sg13g2_decap_8 FILLER_15_1796 ();
 sg13g2_decap_8 FILLER_15_1803 ();
 sg13g2_decap_8 FILLER_15_1810 ();
 sg13g2_decap_8 FILLER_15_1817 ();
 sg13g2_decap_8 FILLER_15_1824 ();
 sg13g2_decap_8 FILLER_15_1831 ();
 sg13g2_decap_8 FILLER_15_1838 ();
 sg13g2_decap_8 FILLER_15_1845 ();
 sg13g2_decap_8 FILLER_15_1852 ();
 sg13g2_decap_8 FILLER_15_1859 ();
 sg13g2_decap_8 FILLER_15_1866 ();
 sg13g2_decap_8 FILLER_15_1873 ();
 sg13g2_decap_8 FILLER_15_1880 ();
 sg13g2_decap_8 FILLER_15_1887 ();
 sg13g2_decap_8 FILLER_15_1894 ();
 sg13g2_decap_8 FILLER_15_1901 ();
 sg13g2_decap_8 FILLER_15_1908 ();
 sg13g2_decap_8 FILLER_15_1915 ();
 sg13g2_decap_8 FILLER_15_1922 ();
 sg13g2_fill_1 FILLER_15_1929 ();
 sg13g2_decap_8 FILLER_15_1955 ();
 sg13g2_decap_8 FILLER_15_1962 ();
 sg13g2_decap_8 FILLER_15_1969 ();
 sg13g2_decap_8 FILLER_15_1976 ();
 sg13g2_fill_2 FILLER_15_1983 ();
 sg13g2_fill_1 FILLER_15_1985 ();
 sg13g2_decap_8 FILLER_15_2011 ();
 sg13g2_decap_8 FILLER_15_2018 ();
 sg13g2_decap_8 FILLER_15_2025 ();
 sg13g2_decap_8 FILLER_15_2032 ();
 sg13g2_decap_8 FILLER_15_2039 ();
 sg13g2_decap_8 FILLER_15_2046 ();
 sg13g2_decap_8 FILLER_15_2053 ();
 sg13g2_decap_8 FILLER_15_2060 ();
 sg13g2_decap_8 FILLER_15_2067 ();
 sg13g2_decap_8 FILLER_15_2074 ();
 sg13g2_decap_8 FILLER_15_2081 ();
 sg13g2_decap_4 FILLER_15_2088 ();
 sg13g2_fill_1 FILLER_15_2092 ();
 sg13g2_decap_8 FILLER_15_2096 ();
 sg13g2_decap_4 FILLER_15_2103 ();
 sg13g2_fill_2 FILLER_15_2107 ();
 sg13g2_decap_8 FILLER_15_2112 ();
 sg13g2_decap_8 FILLER_15_2119 ();
 sg13g2_decap_4 FILLER_15_2126 ();
 sg13g2_fill_2 FILLER_15_2130 ();
 sg13g2_decap_8 FILLER_15_2135 ();
 sg13g2_fill_2 FILLER_15_2142 ();
 sg13g2_fill_1 FILLER_15_2144 ();
 sg13g2_fill_2 FILLER_15_2148 ();
 sg13g2_fill_1 FILLER_15_2150 ();
 sg13g2_decap_8 FILLER_15_2154 ();
 sg13g2_decap_4 FILLER_15_2161 ();
 sg13g2_fill_2 FILLER_15_2165 ();
 sg13g2_decap_8 FILLER_15_2170 ();
 sg13g2_decap_4 FILLER_15_2177 ();
 sg13g2_decap_8 FILLER_15_2184 ();
 sg13g2_decap_8 FILLER_15_2191 ();
 sg13g2_decap_8 FILLER_15_2198 ();
 sg13g2_decap_4 FILLER_15_2205 ();
 sg13g2_fill_1 FILLER_15_2209 ();
 sg13g2_decap_8 FILLER_15_2213 ();
 sg13g2_decap_8 FILLER_15_2220 ();
 sg13g2_decap_8 FILLER_15_2227 ();
 sg13g2_decap_8 FILLER_15_2234 ();
 sg13g2_decap_4 FILLER_15_2241 ();
 sg13g2_fill_1 FILLER_15_2245 ();
 sg13g2_fill_2 FILLER_15_2251 ();
 sg13g2_fill_1 FILLER_15_2253 ();
 sg13g2_decap_8 FILLER_15_2267 ();
 sg13g2_decap_8 FILLER_15_2274 ();
 sg13g2_fill_1 FILLER_15_2281 ();
 sg13g2_fill_2 FILLER_15_2297 ();
 sg13g2_decap_8 FILLER_15_2314 ();
 sg13g2_decap_8 FILLER_15_2321 ();
 sg13g2_decap_8 FILLER_15_2328 ();
 sg13g2_decap_4 FILLER_15_2335 ();
 sg13g2_fill_1 FILLER_15_2339 ();
 sg13g2_decap_4 FILLER_15_2350 ();
 sg13g2_fill_2 FILLER_15_2354 ();
 sg13g2_decap_8 FILLER_15_2360 ();
 sg13g2_fill_2 FILLER_15_2367 ();
 sg13g2_decap_8 FILLER_15_2379 ();
 sg13g2_decap_4 FILLER_15_2386 ();
 sg13g2_decap_4 FILLER_15_2395 ();
 sg13g2_fill_2 FILLER_15_2399 ();
 sg13g2_decap_8 FILLER_15_2414 ();
 sg13g2_decap_4 FILLER_15_2421 ();
 sg13g2_fill_2 FILLER_15_2438 ();
 sg13g2_decap_4 FILLER_15_2466 ();
 sg13g2_fill_1 FILLER_15_2470 ();
 sg13g2_decap_8 FILLER_15_2496 ();
 sg13g2_decap_8 FILLER_15_2528 ();
 sg13g2_decap_8 FILLER_15_2535 ();
 sg13g2_decap_8 FILLER_15_2542 ();
 sg13g2_decap_8 FILLER_15_2549 ();
 sg13g2_decap_8 FILLER_15_2556 ();
 sg13g2_decap_8 FILLER_15_2563 ();
 sg13g2_decap_8 FILLER_15_2570 ();
 sg13g2_decap_8 FILLER_15_2577 ();
 sg13g2_decap_8 FILLER_15_2584 ();
 sg13g2_decap_8 FILLER_15_2591 ();
 sg13g2_decap_8 FILLER_15_2598 ();
 sg13g2_decap_8 FILLER_15_2605 ();
 sg13g2_decap_8 FILLER_15_2612 ();
 sg13g2_decap_8 FILLER_15_2619 ();
 sg13g2_decap_8 FILLER_15_2626 ();
 sg13g2_decap_8 FILLER_15_2633 ();
 sg13g2_decap_8 FILLER_15_2640 ();
 sg13g2_decap_8 FILLER_15_2647 ();
 sg13g2_decap_8 FILLER_15_2654 ();
 sg13g2_decap_8 FILLER_15_2661 ();
 sg13g2_decap_8 FILLER_15_2668 ();
 sg13g2_decap_4 FILLER_15_2675 ();
 sg13g2_decap_8 FILLER_15_2690 ();
 sg13g2_fill_2 FILLER_15_2697 ();
 sg13g2_fill_1 FILLER_15_2699 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_76 ();
 sg13g2_decap_8 FILLER_16_83 ();
 sg13g2_decap_8 FILLER_16_90 ();
 sg13g2_decap_8 FILLER_16_97 ();
 sg13g2_decap_8 FILLER_16_104 ();
 sg13g2_decap_8 FILLER_16_111 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_decap_8 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_decap_8 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_188 ();
 sg13g2_decap_8 FILLER_16_195 ();
 sg13g2_decap_8 FILLER_16_202 ();
 sg13g2_decap_8 FILLER_16_209 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_288 ();
 sg13g2_fill_2 FILLER_16_296 ();
 sg13g2_fill_2 FILLER_16_304 ();
 sg13g2_fill_2 FILLER_16_312 ();
 sg13g2_fill_2 FILLER_16_320 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_344 ();
 sg13g2_fill_2 FILLER_16_352 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_368 ();
 sg13g2_fill_2 FILLER_16_376 ();
 sg13g2_fill_2 FILLER_16_384 ();
 sg13g2_fill_2 FILLER_16_392 ();
 sg13g2_fill_2 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_421 ();
 sg13g2_decap_8 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_16_435 ();
 sg13g2_decap_8 FILLER_16_442 ();
 sg13g2_decap_8 FILLER_16_449 ();
 sg13g2_decap_8 FILLER_16_456 ();
 sg13g2_decap_8 FILLER_16_463 ();
 sg13g2_decap_8 FILLER_16_470 ();
 sg13g2_decap_8 FILLER_16_477 ();
 sg13g2_decap_8 FILLER_16_484 ();
 sg13g2_decap_8 FILLER_16_491 ();
 sg13g2_decap_8 FILLER_16_498 ();
 sg13g2_decap_8 FILLER_16_505 ();
 sg13g2_decap_8 FILLER_16_512 ();
 sg13g2_fill_2 FILLER_16_519 ();
 sg13g2_fill_2 FILLER_16_528 ();
 sg13g2_fill_1 FILLER_16_530 ();
 sg13g2_fill_1 FILLER_16_534 ();
 sg13g2_fill_2 FILLER_16_538 ();
 sg13g2_fill_1 FILLER_16_540 ();
 sg13g2_fill_2 FILLER_16_550 ();
 sg13g2_fill_1 FILLER_16_552 ();
 sg13g2_decap_4 FILLER_16_562 ();
 sg13g2_fill_2 FILLER_16_572 ();
 sg13g2_fill_1 FILLER_16_574 ();
 sg13g2_decap_4 FILLER_16_581 ();
 sg13g2_fill_1 FILLER_16_585 ();
 sg13g2_fill_2 FILLER_16_589 ();
 sg13g2_decap_4 FILLER_16_606 ();
 sg13g2_fill_1 FILLER_16_613 ();
 sg13g2_fill_2 FILLER_16_620 ();
 sg13g2_fill_1 FILLER_16_622 ();
 sg13g2_fill_1 FILLER_16_629 ();
 sg13g2_fill_2 FILLER_16_636 ();
 sg13g2_fill_1 FILLER_16_638 ();
 sg13g2_fill_2 FILLER_16_645 ();
 sg13g2_decap_8 FILLER_16_653 ();
 sg13g2_fill_1 FILLER_16_660 ();
 sg13g2_fill_2 FILLER_16_667 ();
 sg13g2_fill_1 FILLER_16_669 ();
 sg13g2_fill_2 FILLER_16_676 ();
 sg13g2_fill_1 FILLER_16_687 ();
 sg13g2_fill_1 FILLER_16_691 ();
 sg13g2_fill_2 FILLER_16_698 ();
 sg13g2_fill_2 FILLER_16_703 ();
 sg13g2_fill_1 FILLER_16_705 ();
 sg13g2_fill_2 FILLER_16_709 ();
 sg13g2_fill_1 FILLER_16_711 ();
 sg13g2_decap_4 FILLER_16_728 ();
 sg13g2_fill_2 FILLER_16_738 ();
 sg13g2_fill_2 FILLER_16_746 ();
 sg13g2_fill_2 FILLER_16_754 ();
 sg13g2_fill_1 FILLER_16_762 ();
 sg13g2_fill_2 FILLER_16_769 ();
 sg13g2_fill_2 FILLER_16_777 ();
 sg13g2_fill_2 FILLER_16_785 ();
 sg13g2_fill_2 FILLER_16_793 ();
 sg13g2_fill_2 FILLER_16_801 ();
 sg13g2_fill_2 FILLER_16_809 ();
 sg13g2_fill_2 FILLER_16_817 ();
 sg13g2_fill_2 FILLER_16_825 ();
 sg13g2_fill_2 FILLER_16_833 ();
 sg13g2_fill_1 FILLER_16_841 ();
 sg13g2_fill_2 FILLER_16_848 ();
 sg13g2_fill_2 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_864 ();
 sg13g2_fill_1 FILLER_16_866 ();
 sg13g2_decap_8 FILLER_16_872 ();
 sg13g2_decap_8 FILLER_16_879 ();
 sg13g2_decap_8 FILLER_16_886 ();
 sg13g2_decap_8 FILLER_16_893 ();
 sg13g2_decap_8 FILLER_16_900 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_8 FILLER_16_914 ();
 sg13g2_decap_8 FILLER_16_921 ();
 sg13g2_decap_8 FILLER_16_928 ();
 sg13g2_decap_8 FILLER_16_935 ();
 sg13g2_decap_8 FILLER_16_942 ();
 sg13g2_decap_8 FILLER_16_949 ();
 sg13g2_decap_8 FILLER_16_956 ();
 sg13g2_decap_8 FILLER_16_963 ();
 sg13g2_decap_8 FILLER_16_970 ();
 sg13g2_fill_1 FILLER_16_977 ();
 sg13g2_decap_8 FILLER_16_982 ();
 sg13g2_decap_8 FILLER_16_989 ();
 sg13g2_decap_4 FILLER_16_996 ();
 sg13g2_fill_2 FILLER_16_1000 ();
 sg13g2_fill_2 FILLER_16_1008 ();
 sg13g2_fill_1 FILLER_16_1010 ();
 sg13g2_fill_2 FILLER_16_1014 ();
 sg13g2_fill_1 FILLER_16_1019 ();
 sg13g2_decap_8 FILLER_16_1023 ();
 sg13g2_fill_2 FILLER_16_1030 ();
 sg13g2_decap_8 FILLER_16_1035 ();
 sg13g2_decap_4 FILLER_16_1042 ();
 sg13g2_fill_2 FILLER_16_1049 ();
 sg13g2_decap_8 FILLER_16_1054 ();
 sg13g2_fill_1 FILLER_16_1061 ();
 sg13g2_decap_8 FILLER_16_1065 ();
 sg13g2_fill_2 FILLER_16_1072 ();
 sg13g2_fill_1 FILLER_16_1074 ();
 sg13g2_fill_1 FILLER_16_1078 ();
 sg13g2_decap_8 FILLER_16_1082 ();
 sg13g2_decap_8 FILLER_16_1089 ();
 sg13g2_decap_4 FILLER_16_1099 ();
 sg13g2_decap_8 FILLER_16_1106 ();
 sg13g2_decap_4 FILLER_16_1113 ();
 sg13g2_decap_8 FILLER_16_1133 ();
 sg13g2_decap_8 FILLER_16_1140 ();
 sg13g2_decap_8 FILLER_16_1147 ();
 sg13g2_fill_2 FILLER_16_1154 ();
 sg13g2_fill_1 FILLER_16_1156 ();
 sg13g2_fill_2 FILLER_16_1160 ();
 sg13g2_decap_8 FILLER_16_1168 ();
 sg13g2_fill_2 FILLER_16_1181 ();
 sg13g2_fill_2 FILLER_16_1189 ();
 sg13g2_fill_2 FILLER_16_1197 ();
 sg13g2_fill_2 FILLER_16_1205 ();
 sg13g2_fill_2 FILLER_16_1213 ();
 sg13g2_fill_2 FILLER_16_1221 ();
 sg13g2_fill_2 FILLER_16_1229 ();
 sg13g2_fill_2 FILLER_16_1237 ();
 sg13g2_fill_1 FILLER_16_1239 ();
 sg13g2_fill_2 FILLER_16_1246 ();
 sg13g2_fill_2 FILLER_16_1254 ();
 sg13g2_fill_2 FILLER_16_1262 ();
 sg13g2_fill_2 FILLER_16_1270 ();
 sg13g2_fill_2 FILLER_16_1278 ();
 sg13g2_fill_2 FILLER_16_1286 ();
 sg13g2_fill_1 FILLER_16_1306 ();
 sg13g2_fill_2 FILLER_16_1313 ();
 sg13g2_fill_1 FILLER_16_1315 ();
 sg13g2_fill_2 FILLER_16_1322 ();
 sg13g2_decap_8 FILLER_16_1329 ();
 sg13g2_decap_8 FILLER_16_1336 ();
 sg13g2_decap_4 FILLER_16_1343 ();
 sg13g2_decap_8 FILLER_16_1350 ();
 sg13g2_decap_8 FILLER_16_1357 ();
 sg13g2_decap_8 FILLER_16_1364 ();
 sg13g2_fill_2 FILLER_16_1371 ();
 sg13g2_decap_8 FILLER_16_1376 ();
 sg13g2_decap_8 FILLER_16_1383 ();
 sg13g2_decap_8 FILLER_16_1390 ();
 sg13g2_decap_8 FILLER_16_1397 ();
 sg13g2_decap_8 FILLER_16_1404 ();
 sg13g2_decap_8 FILLER_16_1411 ();
 sg13g2_decap_8 FILLER_16_1418 ();
 sg13g2_fill_2 FILLER_16_1425 ();
 sg13g2_decap_8 FILLER_16_1434 ();
 sg13g2_fill_2 FILLER_16_1441 ();
 sg13g2_fill_1 FILLER_16_1443 ();
 sg13g2_decap_4 FILLER_16_1447 ();
 sg13g2_fill_2 FILLER_16_1451 ();
 sg13g2_decap_4 FILLER_16_1456 ();
 sg13g2_fill_1 FILLER_16_1460 ();
 sg13g2_decap_4 FILLER_16_1464 ();
 sg13g2_fill_1 FILLER_16_1468 ();
 sg13g2_decap_8 FILLER_16_1472 ();
 sg13g2_decap_8 FILLER_16_1479 ();
 sg13g2_decap_8 FILLER_16_1486 ();
 sg13g2_decap_8 FILLER_16_1493 ();
 sg13g2_fill_1 FILLER_16_1500 ();
 sg13g2_decap_8 FILLER_16_1504 ();
 sg13g2_decap_4 FILLER_16_1511 ();
 sg13g2_fill_2 FILLER_16_1515 ();
 sg13g2_decap_4 FILLER_16_1520 ();
 sg13g2_fill_1 FILLER_16_1524 ();
 sg13g2_decap_4 FILLER_16_1528 ();
 sg13g2_fill_1 FILLER_16_1532 ();
 sg13g2_decap_4 FILLER_16_1536 ();
 sg13g2_fill_2 FILLER_16_1540 ();
 sg13g2_decap_4 FILLER_16_1545 ();
 sg13g2_fill_2 FILLER_16_1549 ();
 sg13g2_decap_8 FILLER_16_1554 ();
 sg13g2_decap_4 FILLER_16_1561 ();
 sg13g2_fill_1 FILLER_16_1565 ();
 sg13g2_decap_8 FILLER_16_1569 ();
 sg13g2_decap_8 FILLER_16_1576 ();
 sg13g2_decap_4 FILLER_16_1583 ();
 sg13g2_fill_2 FILLER_16_1587 ();
 sg13g2_decap_8 FILLER_16_1592 ();
 sg13g2_decap_8 FILLER_16_1599 ();
 sg13g2_decap_8 FILLER_16_1606 ();
 sg13g2_decap_4 FILLER_16_1613 ();
 sg13g2_fill_2 FILLER_16_1617 ();
 sg13g2_fill_1 FILLER_16_1644 ();
 sg13g2_fill_2 FILLER_16_1651 ();
 sg13g2_fill_2 FILLER_16_1659 ();
 sg13g2_fill_1 FILLER_16_1667 ();
 sg13g2_fill_2 FILLER_16_1674 ();
 sg13g2_fill_2 FILLER_16_1682 ();
 sg13g2_fill_2 FILLER_16_1690 ();
 sg13g2_fill_1 FILLER_16_1692 ();
 sg13g2_fill_2 FILLER_16_1699 ();
 sg13g2_fill_2 FILLER_16_1707 ();
 sg13g2_fill_2 FILLER_16_1715 ();
 sg13g2_fill_2 FILLER_16_1723 ();
 sg13g2_fill_2 FILLER_16_1731 ();
 sg13g2_fill_2 FILLER_16_1739 ();
 sg13g2_fill_2 FILLER_16_1747 ();
 sg13g2_fill_2 FILLER_16_1755 ();
 sg13g2_fill_1 FILLER_16_1763 ();
 sg13g2_decap_8 FILLER_16_1775 ();
 sg13g2_decap_8 FILLER_16_1782 ();
 sg13g2_decap_8 FILLER_16_1789 ();
 sg13g2_decap_8 FILLER_16_1796 ();
 sg13g2_decap_4 FILLER_16_1803 ();
 sg13g2_decap_8 FILLER_16_1820 ();
 sg13g2_decap_8 FILLER_16_1827 ();
 sg13g2_decap_8 FILLER_16_1834 ();
 sg13g2_decap_8 FILLER_16_1841 ();
 sg13g2_decap_8 FILLER_16_1848 ();
 sg13g2_decap_8 FILLER_16_1855 ();
 sg13g2_decap_8 FILLER_16_1862 ();
 sg13g2_decap_8 FILLER_16_1869 ();
 sg13g2_decap_8 FILLER_16_1876 ();
 sg13g2_decap_8 FILLER_16_1887 ();
 sg13g2_decap_8 FILLER_16_1894 ();
 sg13g2_decap_4 FILLER_16_1901 ();
 sg13g2_decap_8 FILLER_16_1911 ();
 sg13g2_decap_8 FILLER_16_1921 ();
 sg13g2_decap_4 FILLER_16_1931 ();
 sg13g2_fill_1 FILLER_16_1935 ();
 sg13g2_decap_8 FILLER_16_1939 ();
 sg13g2_decap_8 FILLER_16_1946 ();
 sg13g2_decap_4 FILLER_16_1953 ();
 sg13g2_fill_2 FILLER_16_1957 ();
 sg13g2_decap_4 FILLER_16_1962 ();
 sg13g2_fill_2 FILLER_16_1978 ();
 sg13g2_decap_4 FILLER_16_1983 ();
 sg13g2_decap_8 FILLER_16_1990 ();
 sg13g2_decap_8 FILLER_16_1997 ();
 sg13g2_decap_4 FILLER_16_2004 ();
 sg13g2_fill_1 FILLER_16_2008 ();
 sg13g2_fill_2 FILLER_16_2015 ();
 sg13g2_decap_4 FILLER_16_2020 ();
 sg13g2_fill_1 FILLER_16_2024 ();
 sg13g2_fill_1 FILLER_16_2028 ();
 sg13g2_fill_2 FILLER_16_2035 ();
 sg13g2_fill_1 FILLER_16_2037 ();
 sg13g2_decap_8 FILLER_16_2041 ();
 sg13g2_decap_8 FILLER_16_2048 ();
 sg13g2_decap_8 FILLER_16_2055 ();
 sg13g2_fill_2 FILLER_16_2068 ();
 sg13g2_fill_1 FILLER_16_2070 ();
 sg13g2_decap_4 FILLER_16_2077 ();
 sg13g2_fill_1 FILLER_16_2081 ();
 sg13g2_fill_2 FILLER_16_2088 ();
 sg13g2_fill_2 FILLER_16_2096 ();
 sg13g2_fill_2 FILLER_16_2104 ();
 sg13g2_fill_1 FILLER_16_2112 ();
 sg13g2_fill_2 FILLER_16_2119 ();
 sg13g2_fill_2 FILLER_16_2127 ();
 sg13g2_fill_2 FILLER_16_2144 ();
 sg13g2_fill_2 FILLER_16_2152 ();
 sg13g2_fill_2 FILLER_16_2160 ();
 sg13g2_fill_2 FILLER_16_2168 ();
 sg13g2_fill_2 FILLER_16_2176 ();
 sg13g2_fill_1 FILLER_16_2184 ();
 sg13g2_fill_2 FILLER_16_2191 ();
 sg13g2_fill_2 FILLER_16_2199 ();
 sg13g2_fill_1 FILLER_16_2201 ();
 sg13g2_fill_1 FILLER_16_2211 ();
 sg13g2_fill_2 FILLER_16_2218 ();
 sg13g2_decap_8 FILLER_16_2231 ();
 sg13g2_decap_8 FILLER_16_2238 ();
 sg13g2_decap_8 FILLER_16_2245 ();
 sg13g2_decap_8 FILLER_16_2252 ();
 sg13g2_fill_2 FILLER_16_2259 ();
 sg13g2_decap_8 FILLER_16_2274 ();
 sg13g2_decap_8 FILLER_16_2281 ();
 sg13g2_decap_8 FILLER_16_2288 ();
 sg13g2_fill_2 FILLER_16_2295 ();
 sg13g2_fill_1 FILLER_16_2297 ();
 sg13g2_decap_8 FILLER_16_2302 ();
 sg13g2_decap_8 FILLER_16_2309 ();
 sg13g2_decap_8 FILLER_16_2316 ();
 sg13g2_decap_8 FILLER_16_2323 ();
 sg13g2_fill_2 FILLER_16_2340 ();
 sg13g2_fill_1 FILLER_16_2342 ();
 sg13g2_decap_4 FILLER_16_2346 ();
 sg13g2_fill_1 FILLER_16_2350 ();
 sg13g2_decap_4 FILLER_16_2354 ();
 sg13g2_fill_1 FILLER_16_2358 ();
 sg13g2_decap_4 FILLER_16_2362 ();
 sg13g2_fill_2 FILLER_16_2366 ();
 sg13g2_fill_2 FILLER_16_2371 ();
 sg13g2_fill_1 FILLER_16_2376 ();
 sg13g2_decap_4 FILLER_16_2380 ();
 sg13g2_fill_2 FILLER_16_2384 ();
 sg13g2_decap_8 FILLER_16_2398 ();
 sg13g2_decap_8 FILLER_16_2405 ();
 sg13g2_decap_8 FILLER_16_2412 ();
 sg13g2_decap_8 FILLER_16_2419 ();
 sg13g2_decap_8 FILLER_16_2426 ();
 sg13g2_decap_8 FILLER_16_2433 ();
 sg13g2_decap_4 FILLER_16_2440 ();
 sg13g2_fill_2 FILLER_16_2444 ();
 sg13g2_decap_8 FILLER_16_2451 ();
 sg13g2_decap_8 FILLER_16_2458 ();
 sg13g2_decap_8 FILLER_16_2465 ();
 sg13g2_decap_8 FILLER_16_2472 ();
 sg13g2_fill_2 FILLER_16_2479 ();
 sg13g2_fill_1 FILLER_16_2481 ();
 sg13g2_decap_8 FILLER_16_2485 ();
 sg13g2_decap_8 FILLER_16_2492 ();
 sg13g2_decap_8 FILLER_16_2499 ();
 sg13g2_decap_8 FILLER_16_2506 ();
 sg13g2_decap_8 FILLER_16_2513 ();
 sg13g2_decap_8 FILLER_16_2520 ();
 sg13g2_decap_4 FILLER_16_2527 ();
 sg13g2_fill_2 FILLER_16_2531 ();
 sg13g2_fill_2 FILLER_16_2539 ();
 sg13g2_fill_1 FILLER_16_2541 ();
 sg13g2_fill_1 FILLER_16_2548 ();
 sg13g2_fill_2 FILLER_16_2555 ();
 sg13g2_decap_4 FILLER_16_2569 ();
 sg13g2_fill_2 FILLER_16_2585 ();
 sg13g2_fill_2 FILLER_16_2593 ();
 sg13g2_fill_1 FILLER_16_2595 ();
 sg13g2_fill_2 FILLER_16_2608 ();
 sg13g2_fill_2 FILLER_16_2616 ();
 sg13g2_fill_1 FILLER_16_2618 ();
 sg13g2_fill_2 FILLER_16_2631 ();
 sg13g2_decap_4 FILLER_16_2645 ();
 sg13g2_fill_1 FILLER_16_2649 ();
 sg13g2_fill_2 FILLER_16_2656 ();
 sg13g2_fill_1 FILLER_16_2658 ();
 sg13g2_decap_8 FILLER_16_2676 ();
 sg13g2_decap_8 FILLER_16_2683 ();
 sg13g2_decap_8 FILLER_16_2690 ();
 sg13g2_fill_2 FILLER_16_2697 ();
 sg13g2_fill_1 FILLER_16_2699 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_8 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_980 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_decap_8 FILLER_17_1029 ();
 sg13g2_decap_8 FILLER_17_1036 ();
 sg13g2_decap_8 FILLER_17_1043 ();
 sg13g2_decap_8 FILLER_17_1050 ();
 sg13g2_decap_8 FILLER_17_1057 ();
 sg13g2_decap_8 FILLER_17_1064 ();
 sg13g2_decap_8 FILLER_17_1071 ();
 sg13g2_decap_8 FILLER_17_1078 ();
 sg13g2_decap_8 FILLER_17_1085 ();
 sg13g2_decap_8 FILLER_17_1092 ();
 sg13g2_decap_8 FILLER_17_1099 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_decap_8 FILLER_17_1120 ();
 sg13g2_decap_8 FILLER_17_1127 ();
 sg13g2_decap_8 FILLER_17_1134 ();
 sg13g2_decap_8 FILLER_17_1141 ();
 sg13g2_decap_8 FILLER_17_1148 ();
 sg13g2_decap_8 FILLER_17_1155 ();
 sg13g2_decap_8 FILLER_17_1162 ();
 sg13g2_decap_8 FILLER_17_1169 ();
 sg13g2_decap_8 FILLER_17_1176 ();
 sg13g2_decap_8 FILLER_17_1183 ();
 sg13g2_decap_8 FILLER_17_1190 ();
 sg13g2_decap_8 FILLER_17_1197 ();
 sg13g2_decap_8 FILLER_17_1204 ();
 sg13g2_decap_8 FILLER_17_1211 ();
 sg13g2_decap_8 FILLER_17_1218 ();
 sg13g2_decap_8 FILLER_17_1225 ();
 sg13g2_decap_8 FILLER_17_1232 ();
 sg13g2_decap_8 FILLER_17_1239 ();
 sg13g2_decap_8 FILLER_17_1246 ();
 sg13g2_decap_8 FILLER_17_1253 ();
 sg13g2_decap_8 FILLER_17_1260 ();
 sg13g2_decap_8 FILLER_17_1267 ();
 sg13g2_decap_8 FILLER_17_1274 ();
 sg13g2_decap_8 FILLER_17_1281 ();
 sg13g2_decap_8 FILLER_17_1288 ();
 sg13g2_decap_8 FILLER_17_1295 ();
 sg13g2_decap_8 FILLER_17_1302 ();
 sg13g2_decap_8 FILLER_17_1309 ();
 sg13g2_decap_8 FILLER_17_1316 ();
 sg13g2_decap_8 FILLER_17_1323 ();
 sg13g2_decap_8 FILLER_17_1330 ();
 sg13g2_decap_8 FILLER_17_1337 ();
 sg13g2_decap_8 FILLER_17_1344 ();
 sg13g2_decap_8 FILLER_17_1351 ();
 sg13g2_decap_8 FILLER_17_1358 ();
 sg13g2_decap_8 FILLER_17_1365 ();
 sg13g2_decap_8 FILLER_17_1372 ();
 sg13g2_decap_8 FILLER_17_1379 ();
 sg13g2_decap_8 FILLER_17_1386 ();
 sg13g2_decap_8 FILLER_17_1393 ();
 sg13g2_decap_8 FILLER_17_1400 ();
 sg13g2_decap_8 FILLER_17_1407 ();
 sg13g2_decap_8 FILLER_17_1414 ();
 sg13g2_decap_8 FILLER_17_1421 ();
 sg13g2_decap_8 FILLER_17_1428 ();
 sg13g2_decap_8 FILLER_17_1435 ();
 sg13g2_decap_8 FILLER_17_1442 ();
 sg13g2_decap_8 FILLER_17_1449 ();
 sg13g2_decap_8 FILLER_17_1456 ();
 sg13g2_decap_8 FILLER_17_1463 ();
 sg13g2_decap_8 FILLER_17_1470 ();
 sg13g2_decap_8 FILLER_17_1477 ();
 sg13g2_decap_8 FILLER_17_1484 ();
 sg13g2_decap_8 FILLER_17_1491 ();
 sg13g2_decap_8 FILLER_17_1498 ();
 sg13g2_decap_8 FILLER_17_1505 ();
 sg13g2_decap_8 FILLER_17_1512 ();
 sg13g2_decap_8 FILLER_17_1519 ();
 sg13g2_decap_8 FILLER_17_1526 ();
 sg13g2_decap_8 FILLER_17_1533 ();
 sg13g2_decap_8 FILLER_17_1540 ();
 sg13g2_decap_8 FILLER_17_1547 ();
 sg13g2_decap_8 FILLER_17_1554 ();
 sg13g2_decap_8 FILLER_17_1561 ();
 sg13g2_decap_8 FILLER_17_1568 ();
 sg13g2_decap_8 FILLER_17_1575 ();
 sg13g2_decap_8 FILLER_17_1582 ();
 sg13g2_decap_8 FILLER_17_1589 ();
 sg13g2_decap_8 FILLER_17_1596 ();
 sg13g2_decap_8 FILLER_17_1603 ();
 sg13g2_decap_8 FILLER_17_1610 ();
 sg13g2_decap_8 FILLER_17_1617 ();
 sg13g2_decap_8 FILLER_17_1624 ();
 sg13g2_decap_8 FILLER_17_1631 ();
 sg13g2_decap_8 FILLER_17_1638 ();
 sg13g2_decap_8 FILLER_17_1645 ();
 sg13g2_decap_8 FILLER_17_1652 ();
 sg13g2_decap_8 FILLER_17_1659 ();
 sg13g2_decap_8 FILLER_17_1666 ();
 sg13g2_decap_8 FILLER_17_1673 ();
 sg13g2_decap_8 FILLER_17_1680 ();
 sg13g2_decap_8 FILLER_17_1687 ();
 sg13g2_decap_8 FILLER_17_1694 ();
 sg13g2_decap_8 FILLER_17_1701 ();
 sg13g2_decap_8 FILLER_17_1708 ();
 sg13g2_decap_8 FILLER_17_1715 ();
 sg13g2_decap_8 FILLER_17_1722 ();
 sg13g2_decap_8 FILLER_17_1729 ();
 sg13g2_decap_8 FILLER_17_1736 ();
 sg13g2_decap_8 FILLER_17_1743 ();
 sg13g2_decap_8 FILLER_17_1750 ();
 sg13g2_decap_8 FILLER_17_1757 ();
 sg13g2_decap_8 FILLER_17_1764 ();
 sg13g2_decap_8 FILLER_17_1771 ();
 sg13g2_decap_8 FILLER_17_1778 ();
 sg13g2_decap_8 FILLER_17_1785 ();
 sg13g2_decap_8 FILLER_17_1792 ();
 sg13g2_decap_8 FILLER_17_1799 ();
 sg13g2_decap_8 FILLER_17_1806 ();
 sg13g2_decap_8 FILLER_17_1813 ();
 sg13g2_decap_8 FILLER_17_1820 ();
 sg13g2_decap_8 FILLER_17_1827 ();
 sg13g2_decap_8 FILLER_17_1834 ();
 sg13g2_decap_8 FILLER_17_1841 ();
 sg13g2_decap_8 FILLER_17_1848 ();
 sg13g2_decap_8 FILLER_17_1855 ();
 sg13g2_decap_8 FILLER_17_1862 ();
 sg13g2_decap_8 FILLER_17_1869 ();
 sg13g2_decap_8 FILLER_17_1876 ();
 sg13g2_decap_8 FILLER_17_1883 ();
 sg13g2_decap_8 FILLER_17_1890 ();
 sg13g2_decap_8 FILLER_17_1897 ();
 sg13g2_decap_8 FILLER_17_1904 ();
 sg13g2_decap_8 FILLER_17_1911 ();
 sg13g2_decap_8 FILLER_17_1918 ();
 sg13g2_decap_8 FILLER_17_1925 ();
 sg13g2_decap_8 FILLER_17_1932 ();
 sg13g2_decap_8 FILLER_17_1939 ();
 sg13g2_decap_8 FILLER_17_1946 ();
 sg13g2_decap_8 FILLER_17_1953 ();
 sg13g2_decap_8 FILLER_17_1960 ();
 sg13g2_decap_8 FILLER_17_1967 ();
 sg13g2_decap_8 FILLER_17_1974 ();
 sg13g2_decap_8 FILLER_17_1981 ();
 sg13g2_decap_8 FILLER_17_1988 ();
 sg13g2_decap_8 FILLER_17_1995 ();
 sg13g2_decap_8 FILLER_17_2002 ();
 sg13g2_decap_8 FILLER_17_2009 ();
 sg13g2_decap_8 FILLER_17_2016 ();
 sg13g2_decap_8 FILLER_17_2023 ();
 sg13g2_decap_8 FILLER_17_2030 ();
 sg13g2_decap_8 FILLER_17_2037 ();
 sg13g2_decap_8 FILLER_17_2044 ();
 sg13g2_decap_8 FILLER_17_2051 ();
 sg13g2_decap_8 FILLER_17_2058 ();
 sg13g2_decap_8 FILLER_17_2065 ();
 sg13g2_decap_8 FILLER_17_2072 ();
 sg13g2_decap_8 FILLER_17_2079 ();
 sg13g2_decap_8 FILLER_17_2086 ();
 sg13g2_fill_2 FILLER_17_2093 ();
 sg13g2_decap_8 FILLER_17_2098 ();
 sg13g2_decap_8 FILLER_17_2105 ();
 sg13g2_decap_8 FILLER_17_2112 ();
 sg13g2_decap_8 FILLER_17_2119 ();
 sg13g2_decap_8 FILLER_17_2126 ();
 sg13g2_decap_8 FILLER_17_2133 ();
 sg13g2_decap_8 FILLER_17_2140 ();
 sg13g2_decap_8 FILLER_17_2147 ();
 sg13g2_decap_8 FILLER_17_2154 ();
 sg13g2_decap_8 FILLER_17_2161 ();
 sg13g2_decap_8 FILLER_17_2168 ();
 sg13g2_decap_8 FILLER_17_2175 ();
 sg13g2_decap_8 FILLER_17_2182 ();
 sg13g2_decap_8 FILLER_17_2189 ();
 sg13g2_decap_8 FILLER_17_2196 ();
 sg13g2_decap_8 FILLER_17_2203 ();
 sg13g2_decap_8 FILLER_17_2210 ();
 sg13g2_decap_8 FILLER_17_2217 ();
 sg13g2_decap_8 FILLER_17_2224 ();
 sg13g2_decap_8 FILLER_17_2231 ();
 sg13g2_decap_8 FILLER_17_2238 ();
 sg13g2_decap_8 FILLER_17_2245 ();
 sg13g2_decap_8 FILLER_17_2252 ();
 sg13g2_decap_8 FILLER_17_2259 ();
 sg13g2_decap_8 FILLER_17_2266 ();
 sg13g2_decap_8 FILLER_17_2273 ();
 sg13g2_decap_8 FILLER_17_2280 ();
 sg13g2_decap_8 FILLER_17_2287 ();
 sg13g2_decap_8 FILLER_17_2294 ();
 sg13g2_decap_8 FILLER_17_2301 ();
 sg13g2_decap_8 FILLER_17_2308 ();
 sg13g2_decap_8 FILLER_17_2315 ();
 sg13g2_decap_8 FILLER_17_2322 ();
 sg13g2_decap_8 FILLER_17_2329 ();
 sg13g2_decap_8 FILLER_17_2336 ();
 sg13g2_decap_8 FILLER_17_2343 ();
 sg13g2_decap_8 FILLER_17_2350 ();
 sg13g2_decap_8 FILLER_17_2357 ();
 sg13g2_decap_8 FILLER_17_2364 ();
 sg13g2_decap_8 FILLER_17_2371 ();
 sg13g2_decap_8 FILLER_17_2378 ();
 sg13g2_decap_8 FILLER_17_2385 ();
 sg13g2_decap_8 FILLER_17_2392 ();
 sg13g2_decap_8 FILLER_17_2399 ();
 sg13g2_decap_8 FILLER_17_2406 ();
 sg13g2_decap_8 FILLER_17_2413 ();
 sg13g2_decap_8 FILLER_17_2420 ();
 sg13g2_decap_8 FILLER_17_2427 ();
 sg13g2_decap_8 FILLER_17_2434 ();
 sg13g2_decap_8 FILLER_17_2441 ();
 sg13g2_decap_8 FILLER_17_2448 ();
 sg13g2_decap_8 FILLER_17_2455 ();
 sg13g2_decap_8 FILLER_17_2462 ();
 sg13g2_decap_8 FILLER_17_2469 ();
 sg13g2_decap_8 FILLER_17_2476 ();
 sg13g2_decap_8 FILLER_17_2483 ();
 sg13g2_decap_8 FILLER_17_2490 ();
 sg13g2_decap_8 FILLER_17_2497 ();
 sg13g2_decap_8 FILLER_17_2504 ();
 sg13g2_decap_8 FILLER_17_2511 ();
 sg13g2_decap_8 FILLER_17_2518 ();
 sg13g2_decap_8 FILLER_17_2525 ();
 sg13g2_decap_8 FILLER_17_2532 ();
 sg13g2_decap_8 FILLER_17_2539 ();
 sg13g2_decap_8 FILLER_17_2546 ();
 sg13g2_decap_8 FILLER_17_2553 ();
 sg13g2_decap_8 FILLER_17_2560 ();
 sg13g2_decap_8 FILLER_17_2567 ();
 sg13g2_decap_8 FILLER_17_2574 ();
 sg13g2_decap_8 FILLER_17_2581 ();
 sg13g2_decap_8 FILLER_17_2588 ();
 sg13g2_decap_8 FILLER_17_2595 ();
 sg13g2_decap_8 FILLER_17_2602 ();
 sg13g2_decap_8 FILLER_17_2609 ();
 sg13g2_decap_8 FILLER_17_2616 ();
 sg13g2_decap_8 FILLER_17_2623 ();
 sg13g2_decap_8 FILLER_17_2630 ();
 sg13g2_decap_8 FILLER_17_2637 ();
 sg13g2_decap_8 FILLER_17_2644 ();
 sg13g2_decap_8 FILLER_17_2651 ();
 sg13g2_decap_8 FILLER_17_2658 ();
 sg13g2_decap_8 FILLER_17_2665 ();
 sg13g2_decap_8 FILLER_17_2672 ();
 sg13g2_decap_8 FILLER_17_2679 ();
 sg13g2_decap_8 FILLER_17_2686 ();
 sg13g2_decap_8 FILLER_17_2693 ();
 assign um_k_zero[0] = \block[0].tie_I.lo ;
 assign um_ena[0] = \block[0].zbuf_ena_I.z ;
 assign um_iw[0] = \block[0].zbuf_iw_I[0].z ;
 assign um_iw[10] = \block[0].zbuf_iw_I[10].z ;
 assign um_iw[11] = \block[0].zbuf_iw_I[11].z ;
 assign um_iw[12] = \block[0].zbuf_iw_I[12].z ;
 assign um_iw[13] = \block[0].zbuf_iw_I[13].z ;
 assign um_iw[14] = \block[0].zbuf_iw_I[14].z ;
 assign um_iw[15] = \block[0].zbuf_iw_I[15].z ;
 assign um_iw[16] = \block[0].zbuf_iw_I[16].z ;
 assign um_iw[17] = \block[0].zbuf_iw_I[17].z ;
 assign um_iw[1] = \block[0].zbuf_iw_I[1].z ;
 assign um_iw[2] = \block[0].zbuf_iw_I[2].z ;
 assign um_iw[3] = \block[0].zbuf_iw_I[3].z ;
 assign um_iw[4] = \block[0].zbuf_iw_I[4].z ;
 assign um_iw[5] = \block[0].zbuf_iw_I[5].z ;
 assign um_iw[6] = \block[0].zbuf_iw_I[6].z ;
 assign um_iw[7] = \block[0].zbuf_iw_I[7].z ;
 assign um_iw[8] = \block[0].zbuf_iw_I[8].z ;
 assign um_iw[9] = \block[0].zbuf_iw_I[9].z ;
 assign um_pg_ena[0] = \block[0].zbuf_pg_ena_I.z ;
 assign um_k_zero[10] = \block[10].tie_I.lo ;
 assign um_ena[10] = \block[10].zbuf_ena_I.z ;
 assign um_iw[180] = \block[10].zbuf_iw_I[0].z ;
 assign um_iw[190] = \block[10].zbuf_iw_I[10].z ;
 assign um_iw[191] = \block[10].zbuf_iw_I[11].z ;
 assign um_iw[192] = \block[10].zbuf_iw_I[12].z ;
 assign um_iw[193] = \block[10].zbuf_iw_I[13].z ;
 assign um_iw[194] = \block[10].zbuf_iw_I[14].z ;
 assign um_iw[195] = \block[10].zbuf_iw_I[15].z ;
 assign um_iw[196] = \block[10].zbuf_iw_I[16].z ;
 assign um_iw[197] = \block[10].zbuf_iw_I[17].z ;
 assign um_iw[181] = \block[10].zbuf_iw_I[1].z ;
 assign um_iw[182] = \block[10].zbuf_iw_I[2].z ;
 assign um_iw[183] = \block[10].zbuf_iw_I[3].z ;
 assign um_iw[184] = \block[10].zbuf_iw_I[4].z ;
 assign um_iw[185] = \block[10].zbuf_iw_I[5].z ;
 assign um_iw[186] = \block[10].zbuf_iw_I[6].z ;
 assign um_iw[187] = \block[10].zbuf_iw_I[7].z ;
 assign um_iw[188] = \block[10].zbuf_iw_I[8].z ;
 assign um_iw[189] = \block[10].zbuf_iw_I[9].z ;
 assign um_pg_ena[10] = \block[10].zbuf_pg_ena_I.z ;
 assign um_k_zero[11] = \block[11].tie_I.lo ;
 assign um_ena[11] = \block[11].zbuf_ena_I.z ;
 assign um_iw[198] = \block[11].zbuf_iw_I[0].z ;
 assign um_iw[208] = \block[11].zbuf_iw_I[10].z ;
 assign um_iw[209] = \block[11].zbuf_iw_I[11].z ;
 assign um_iw[210] = \block[11].zbuf_iw_I[12].z ;
 assign um_iw[211] = \block[11].zbuf_iw_I[13].z ;
 assign um_iw[212] = \block[11].zbuf_iw_I[14].z ;
 assign um_iw[213] = \block[11].zbuf_iw_I[15].z ;
 assign um_iw[214] = \block[11].zbuf_iw_I[16].z ;
 assign um_iw[215] = \block[11].zbuf_iw_I[17].z ;
 assign um_iw[199] = \block[11].zbuf_iw_I[1].z ;
 assign um_iw[200] = \block[11].zbuf_iw_I[2].z ;
 assign um_iw[201] = \block[11].zbuf_iw_I[3].z ;
 assign um_iw[202] = \block[11].zbuf_iw_I[4].z ;
 assign um_iw[203] = \block[11].zbuf_iw_I[5].z ;
 assign um_iw[204] = \block[11].zbuf_iw_I[6].z ;
 assign um_iw[205] = \block[11].zbuf_iw_I[7].z ;
 assign um_iw[206] = \block[11].zbuf_iw_I[8].z ;
 assign um_iw[207] = \block[11].zbuf_iw_I[9].z ;
 assign um_pg_ena[11] = \block[11].zbuf_pg_ena_I.z ;
 assign um_k_zero[1] = \block[1].tie_I.lo ;
 assign um_ena[1] = \block[1].zbuf_ena_I.z ;
 assign um_iw[18] = \block[1].zbuf_iw_I[0].z ;
 assign um_iw[28] = \block[1].zbuf_iw_I[10].z ;
 assign um_iw[29] = \block[1].zbuf_iw_I[11].z ;
 assign um_iw[30] = \block[1].zbuf_iw_I[12].z ;
 assign um_iw[31] = \block[1].zbuf_iw_I[13].z ;
 assign um_iw[32] = \block[1].zbuf_iw_I[14].z ;
 assign um_iw[33] = \block[1].zbuf_iw_I[15].z ;
 assign um_iw[34] = \block[1].zbuf_iw_I[16].z ;
 assign um_iw[35] = \block[1].zbuf_iw_I[17].z ;
 assign um_iw[19] = \block[1].zbuf_iw_I[1].z ;
 assign um_iw[20] = \block[1].zbuf_iw_I[2].z ;
 assign um_iw[21] = \block[1].zbuf_iw_I[3].z ;
 assign um_iw[22] = \block[1].zbuf_iw_I[4].z ;
 assign um_iw[23] = \block[1].zbuf_iw_I[5].z ;
 assign um_iw[24] = \block[1].zbuf_iw_I[6].z ;
 assign um_iw[25] = \block[1].zbuf_iw_I[7].z ;
 assign um_iw[26] = \block[1].zbuf_iw_I[8].z ;
 assign um_iw[27] = \block[1].zbuf_iw_I[9].z ;
 assign um_pg_ena[1] = \block[1].zbuf_pg_ena_I.z ;
 assign um_k_zero[2] = \block[2].tie_I.lo ;
 assign um_ena[2] = \block[2].zbuf_ena_I.z ;
 assign um_iw[36] = \block[2].zbuf_iw_I[0].z ;
 assign um_iw[46] = \block[2].zbuf_iw_I[10].z ;
 assign um_iw[47] = \block[2].zbuf_iw_I[11].z ;
 assign um_iw[48] = \block[2].zbuf_iw_I[12].z ;
 assign um_iw[49] = \block[2].zbuf_iw_I[13].z ;
 assign um_iw[50] = \block[2].zbuf_iw_I[14].z ;
 assign um_iw[51] = \block[2].zbuf_iw_I[15].z ;
 assign um_iw[52] = \block[2].zbuf_iw_I[16].z ;
 assign um_iw[53] = \block[2].zbuf_iw_I[17].z ;
 assign um_iw[37] = \block[2].zbuf_iw_I[1].z ;
 assign um_iw[38] = \block[2].zbuf_iw_I[2].z ;
 assign um_iw[39] = \block[2].zbuf_iw_I[3].z ;
 assign um_iw[40] = \block[2].zbuf_iw_I[4].z ;
 assign um_iw[41] = \block[2].zbuf_iw_I[5].z ;
 assign um_iw[42] = \block[2].zbuf_iw_I[6].z ;
 assign um_iw[43] = \block[2].zbuf_iw_I[7].z ;
 assign um_iw[44] = \block[2].zbuf_iw_I[8].z ;
 assign um_iw[45] = \block[2].zbuf_iw_I[9].z ;
 assign um_pg_ena[2] = \block[2].zbuf_pg_ena_I.z ;
 assign um_k_zero[3] = \block[3].tie_I.lo ;
 assign um_ena[3] = \block[3].zbuf_ena_I.z ;
 assign um_iw[54] = \block[3].zbuf_iw_I[0].z ;
 assign um_iw[64] = \block[3].zbuf_iw_I[10].z ;
 assign um_iw[65] = \block[3].zbuf_iw_I[11].z ;
 assign um_iw[66] = \block[3].zbuf_iw_I[12].z ;
 assign um_iw[67] = \block[3].zbuf_iw_I[13].z ;
 assign um_iw[68] = \block[3].zbuf_iw_I[14].z ;
 assign um_iw[69] = \block[3].zbuf_iw_I[15].z ;
 assign um_iw[70] = \block[3].zbuf_iw_I[16].z ;
 assign um_iw[71] = \block[3].zbuf_iw_I[17].z ;
 assign um_iw[55] = \block[3].zbuf_iw_I[1].z ;
 assign um_iw[56] = \block[3].zbuf_iw_I[2].z ;
 assign um_iw[57] = \block[3].zbuf_iw_I[3].z ;
 assign um_iw[58] = \block[3].zbuf_iw_I[4].z ;
 assign um_iw[59] = \block[3].zbuf_iw_I[5].z ;
 assign um_iw[60] = \block[3].zbuf_iw_I[6].z ;
 assign um_iw[61] = \block[3].zbuf_iw_I[7].z ;
 assign um_iw[62] = \block[3].zbuf_iw_I[8].z ;
 assign um_iw[63] = \block[3].zbuf_iw_I[9].z ;
 assign um_pg_ena[3] = \block[3].zbuf_pg_ena_I.z ;
 assign um_k_zero[4] = \block[4].tie_I.lo ;
 assign um_ena[4] = \block[4].zbuf_ena_I.z ;
 assign um_iw[72] = \block[4].zbuf_iw_I[0].z ;
 assign um_iw[82] = \block[4].zbuf_iw_I[10].z ;
 assign um_iw[83] = \block[4].zbuf_iw_I[11].z ;
 assign um_iw[84] = \block[4].zbuf_iw_I[12].z ;
 assign um_iw[85] = \block[4].zbuf_iw_I[13].z ;
 assign um_iw[86] = \block[4].zbuf_iw_I[14].z ;
 assign um_iw[87] = \block[4].zbuf_iw_I[15].z ;
 assign um_iw[88] = \block[4].zbuf_iw_I[16].z ;
 assign um_iw[89] = \block[4].zbuf_iw_I[17].z ;
 assign um_iw[73] = \block[4].zbuf_iw_I[1].z ;
 assign um_iw[74] = \block[4].zbuf_iw_I[2].z ;
 assign um_iw[75] = \block[4].zbuf_iw_I[3].z ;
 assign um_iw[76] = \block[4].zbuf_iw_I[4].z ;
 assign um_iw[77] = \block[4].zbuf_iw_I[5].z ;
 assign um_iw[78] = \block[4].zbuf_iw_I[6].z ;
 assign um_iw[79] = \block[4].zbuf_iw_I[7].z ;
 assign um_iw[80] = \block[4].zbuf_iw_I[8].z ;
 assign um_iw[81] = \block[4].zbuf_iw_I[9].z ;
 assign um_pg_ena[4] = \block[4].zbuf_pg_ena_I.z ;
 assign um_k_zero[5] = \block[5].tie_I.lo ;
 assign um_ena[5] = \block[5].zbuf_ena_I.z ;
 assign um_iw[90] = \block[5].zbuf_iw_I[0].z ;
 assign um_iw[100] = \block[5].zbuf_iw_I[10].z ;
 assign um_iw[101] = \block[5].zbuf_iw_I[11].z ;
 assign um_iw[102] = \block[5].zbuf_iw_I[12].z ;
 assign um_iw[103] = \block[5].zbuf_iw_I[13].z ;
 assign um_iw[104] = \block[5].zbuf_iw_I[14].z ;
 assign um_iw[105] = \block[5].zbuf_iw_I[15].z ;
 assign um_iw[106] = \block[5].zbuf_iw_I[16].z ;
 assign um_iw[107] = \block[5].zbuf_iw_I[17].z ;
 assign um_iw[91] = \block[5].zbuf_iw_I[1].z ;
 assign um_iw[92] = \block[5].zbuf_iw_I[2].z ;
 assign um_iw[93] = \block[5].zbuf_iw_I[3].z ;
 assign um_iw[94] = \block[5].zbuf_iw_I[4].z ;
 assign um_iw[95] = \block[5].zbuf_iw_I[5].z ;
 assign um_iw[96] = \block[5].zbuf_iw_I[6].z ;
 assign um_iw[97] = \block[5].zbuf_iw_I[7].z ;
 assign um_iw[98] = \block[5].zbuf_iw_I[8].z ;
 assign um_iw[99] = \block[5].zbuf_iw_I[9].z ;
 assign um_pg_ena[5] = \block[5].zbuf_pg_ena_I.z ;
 assign um_k_zero[6] = \block[6].tie_I.lo ;
 assign um_ena[6] = \block[6].zbuf_ena_I.z ;
 assign um_iw[108] = \block[6].zbuf_iw_I[0].z ;
 assign um_iw[118] = \block[6].zbuf_iw_I[10].z ;
 assign um_iw[119] = \block[6].zbuf_iw_I[11].z ;
 assign um_iw[120] = \block[6].zbuf_iw_I[12].z ;
 assign um_iw[121] = \block[6].zbuf_iw_I[13].z ;
 assign um_iw[122] = \block[6].zbuf_iw_I[14].z ;
 assign um_iw[123] = \block[6].zbuf_iw_I[15].z ;
 assign um_iw[124] = \block[6].zbuf_iw_I[16].z ;
 assign um_iw[125] = \block[6].zbuf_iw_I[17].z ;
 assign um_iw[109] = \block[6].zbuf_iw_I[1].z ;
 assign um_iw[110] = \block[6].zbuf_iw_I[2].z ;
 assign um_iw[111] = \block[6].zbuf_iw_I[3].z ;
 assign um_iw[112] = \block[6].zbuf_iw_I[4].z ;
 assign um_iw[113] = \block[6].zbuf_iw_I[5].z ;
 assign um_iw[114] = \block[6].zbuf_iw_I[6].z ;
 assign um_iw[115] = \block[6].zbuf_iw_I[7].z ;
 assign um_iw[116] = \block[6].zbuf_iw_I[8].z ;
 assign um_iw[117] = \block[6].zbuf_iw_I[9].z ;
 assign um_pg_ena[6] = \block[6].zbuf_pg_ena_I.z ;
 assign um_k_zero[7] = \block[7].tie_I.lo ;
 assign um_ena[7] = \block[7].zbuf_ena_I.z ;
 assign um_iw[126] = \block[7].zbuf_iw_I[0].z ;
 assign um_iw[136] = \block[7].zbuf_iw_I[10].z ;
 assign um_iw[137] = \block[7].zbuf_iw_I[11].z ;
 assign um_iw[138] = \block[7].zbuf_iw_I[12].z ;
 assign um_iw[139] = \block[7].zbuf_iw_I[13].z ;
 assign um_iw[140] = \block[7].zbuf_iw_I[14].z ;
 assign um_iw[141] = \block[7].zbuf_iw_I[15].z ;
 assign um_iw[142] = \block[7].zbuf_iw_I[16].z ;
 assign um_iw[143] = \block[7].zbuf_iw_I[17].z ;
 assign um_iw[127] = \block[7].zbuf_iw_I[1].z ;
 assign um_iw[128] = \block[7].zbuf_iw_I[2].z ;
 assign um_iw[129] = \block[7].zbuf_iw_I[3].z ;
 assign um_iw[130] = \block[7].zbuf_iw_I[4].z ;
 assign um_iw[131] = \block[7].zbuf_iw_I[5].z ;
 assign um_iw[132] = \block[7].zbuf_iw_I[6].z ;
 assign um_iw[133] = \block[7].zbuf_iw_I[7].z ;
 assign um_iw[134] = \block[7].zbuf_iw_I[8].z ;
 assign um_iw[135] = \block[7].zbuf_iw_I[9].z ;
 assign um_pg_ena[7] = \block[7].zbuf_pg_ena_I.z ;
 assign um_k_zero[8] = \block[8].tie_I.lo ;
 assign um_ena[8] = \block[8].zbuf_ena_I.z ;
 assign um_iw[144] = \block[8].zbuf_iw_I[0].z ;
 assign um_iw[154] = \block[8].zbuf_iw_I[10].z ;
 assign um_iw[155] = \block[8].zbuf_iw_I[11].z ;
 assign um_iw[156] = \block[8].zbuf_iw_I[12].z ;
 assign um_iw[157] = \block[8].zbuf_iw_I[13].z ;
 assign um_iw[158] = \block[8].zbuf_iw_I[14].z ;
 assign um_iw[159] = \block[8].zbuf_iw_I[15].z ;
 assign um_iw[160] = \block[8].zbuf_iw_I[16].z ;
 assign um_iw[161] = \block[8].zbuf_iw_I[17].z ;
 assign um_iw[145] = \block[8].zbuf_iw_I[1].z ;
 assign um_iw[146] = \block[8].zbuf_iw_I[2].z ;
 assign um_iw[147] = \block[8].zbuf_iw_I[3].z ;
 assign um_iw[148] = \block[8].zbuf_iw_I[4].z ;
 assign um_iw[149] = \block[8].zbuf_iw_I[5].z ;
 assign um_iw[150] = \block[8].zbuf_iw_I[6].z ;
 assign um_iw[151] = \block[8].zbuf_iw_I[7].z ;
 assign um_iw[152] = \block[8].zbuf_iw_I[8].z ;
 assign um_iw[153] = \block[8].zbuf_iw_I[9].z ;
 assign um_pg_ena[8] = \block[8].zbuf_pg_ena_I.z ;
 assign um_k_zero[9] = \block[9].tie_I.lo ;
 assign um_ena[9] = \block[9].zbuf_ena_I.z ;
 assign um_iw[162] = \block[9].zbuf_iw_I[0].z ;
 assign um_iw[172] = \block[9].zbuf_iw_I[10].z ;
 assign um_iw[173] = \block[9].zbuf_iw_I[11].z ;
 assign um_iw[174] = \block[9].zbuf_iw_I[12].z ;
 assign um_iw[175] = \block[9].zbuf_iw_I[13].z ;
 assign um_iw[176] = \block[9].zbuf_iw_I[14].z ;
 assign um_iw[177] = \block[9].zbuf_iw_I[15].z ;
 assign um_iw[178] = \block[9].zbuf_iw_I[16].z ;
 assign um_iw[179] = \block[9].zbuf_iw_I[17].z ;
 assign um_iw[163] = \block[9].zbuf_iw_I[1].z ;
 assign um_iw[164] = \block[9].zbuf_iw_I[2].z ;
 assign um_iw[165] = \block[9].zbuf_iw_I[3].z ;
 assign um_iw[166] = \block[9].zbuf_iw_I[4].z ;
 assign um_iw[167] = \block[9].zbuf_iw_I[5].z ;
 assign um_iw[168] = \block[9].zbuf_iw_I[6].z ;
 assign um_iw[169] = \block[9].zbuf_iw_I[7].z ;
 assign um_iw[170] = \block[9].zbuf_iw_I[8].z ;
 assign um_iw[171] = \block[9].zbuf_iw_I[9].z ;
 assign um_pg_ena[9] = \block[9].zbuf_pg_ena_I.z ;
 assign spine_ow[25] = so_gh;
 assign spine_ow[0] = so_gl;
 assign spine_ow[1] = \tbuf_spine_ow_I[0].z ;
 assign spine_ow[11] = \tbuf_spine_ow_I[10].z ;
 assign spine_ow[12] = \tbuf_spine_ow_I[11].z ;
 assign spine_ow[13] = \tbuf_spine_ow_I[12].z ;
 assign spine_ow[14] = \tbuf_spine_ow_I[13].z ;
 assign spine_ow[15] = \tbuf_spine_ow_I[14].z ;
 assign spine_ow[16] = \tbuf_spine_ow_I[15].z ;
 assign spine_ow[17] = \tbuf_spine_ow_I[16].z ;
 assign spine_ow[18] = \tbuf_spine_ow_I[17].z ;
 assign spine_ow[19] = \tbuf_spine_ow_I[18].z ;
 assign spine_ow[20] = \tbuf_spine_ow_I[19].z ;
 assign spine_ow[2] = \tbuf_spine_ow_I[1].z ;
 assign spine_ow[21] = \tbuf_spine_ow_I[20].z ;
 assign spine_ow[22] = \tbuf_spine_ow_I[21].z ;
 assign spine_ow[23] = \tbuf_spine_ow_I[22].z ;
 assign spine_ow[24] = \tbuf_spine_ow_I[23].z ;
 assign spine_ow[3] = \tbuf_spine_ow_I[2].z ;
 assign spine_ow[4] = \tbuf_spine_ow_I[3].z ;
 assign spine_ow[5] = \tbuf_spine_ow_I[4].z ;
 assign spine_ow[6] = \tbuf_spine_ow_I[5].z ;
 assign spine_ow[7] = \tbuf_spine_ow_I[6].z ;
 assign spine_ow[8] = \tbuf_spine_ow_I[7].z ;
 assign spine_ow[9] = \tbuf_spine_ow_I[8].z ;
 assign spine_ow[10] = \tbuf_spine_ow_I[9].z ;
endmodule
