module tt_ctrl (ctrl_ena,
    ctrl_sel_inc,
    ctrl_sel_rst_n,
    k_one,
    k_zero,
    pad_ui_in,
    pad_uio_in,
    pad_uio_oex,
    pad_uio_out,
    pad_uo_out,
    spine_bot_iw,
    spine_bot_ow,
    spine_top_iw,
    spine_top_ow);
 input ctrl_ena;
 input ctrl_sel_inc;
 input ctrl_sel_rst_n;
 output k_one;
 output k_zero;
 input [9:0] pad_ui_in;
 input [7:0] pad_uio_in;
 output [7:0] pad_uio_oex;
 output [7:0] pad_uio_out;
 output [7:0] pad_uo_out;
 output [29:0] spine_bot_iw;
 input [25:0] spine_bot_ow;
 output [29:0] spine_top_iw;
 input [25:0] spine_top_ow;

 wire ctrl_ena_ibuf;
 wire \ctrl_ibuf_I[1].z ;
 wire \ctrl_ibuf_I[2].z ;
 wire \genblk1[0].pull ;
 wire \genblk1[0].tbuf_pol_spine_ow_I.tx ;
 wire \genblk1[0].tbuf_spine_ow_I[0].a ;
 wire \genblk1[1].pull ;
 wire \genblk1[1].tbuf_pol_spine_ow_I.tx ;
 wire \genblk1[1].tbuf_spine_ow_I[0].a ;
 wire \genblk2[0].ctrl_ena_buf_I.a ;
 wire \genblk2[0].ctrl_ena_buf_I.z ;
 wire \genblk2[0].pad_ui_in_buf_I[0].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[0].z ;
 wire \genblk2[0].pad_ui_in_buf_I[1].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[1].z ;
 wire \genblk2[0].pad_ui_in_buf_I[2].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[2].z ;
 wire \genblk2[0].pad_ui_in_buf_I[3].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[3].z ;
 wire \genblk2[0].pad_ui_in_buf_I[4].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[4].z ;
 wire \genblk2[0].pad_ui_in_buf_I[5].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[5].z ;
 wire \genblk2[0].pad_ui_in_buf_I[6].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[6].z ;
 wire \genblk2[0].pad_ui_in_buf_I[7].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[7].z ;
 wire \genblk2[0].pad_ui_in_buf_I[8].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[8].z ;
 wire \genblk2[0].pad_ui_in_buf_I[9].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[9].z ;
 wire \genblk2[0].pad_uio_in_buf_I[0].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[0].z ;
 wire \genblk2[0].pad_uio_in_buf_I[1].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[1].z ;
 wire \genblk2[0].pad_uio_in_buf_I[2].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[2].z ;
 wire \genblk2[0].pad_uio_in_buf_I[3].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[3].z ;
 wire \genblk2[0].pad_uio_in_buf_I[4].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[4].z ;
 wire \genblk2[0].pad_uio_in_buf_I[5].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[5].z ;
 wire \genblk2[0].pad_uio_in_buf_I[6].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[6].z ;
 wire \genblk2[0].pad_uio_in_buf_I[7].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[7].z ;
 wire \genblk2[0].sel_cnt_buf_I[0].a ;
 wire \genblk2[0].sel_cnt_buf_I[0].z ;
 wire \genblk2[0].sel_cnt_buf_I[1].a ;
 wire \genblk2[0].sel_cnt_buf_I[1].z ;
 wire \genblk2[0].sel_cnt_buf_I[2].a ;
 wire \genblk2[0].sel_cnt_buf_I[2].z ;
 wire \genblk2[0].sel_cnt_buf_I[3].a ;
 wire \genblk2[0].sel_cnt_buf_I[3].z ;
 wire \genblk2[0].sel_cnt_buf_I[4].a ;
 wire \genblk2[0].sel_cnt_buf_I[4].z ;
 wire \genblk2[0].sel_cnt_buf_I[5].a ;
 wire \genblk2[0].sel_cnt_buf_I[5].z ;
 wire \genblk2[0].sel_cnt_buf_I[6].a ;
 wire \genblk2[0].sel_cnt_buf_I[6].z ;
 wire \genblk2[0].sel_cnt_buf_I[7].a ;
 wire \genblk2[0].sel_cnt_buf_I[7].z ;
 wire \genblk2[0].sel_cnt_buf_I[8].a ;
 wire \genblk2[0].sel_cnt_buf_I[8].z ;
 wire \genblk2[0].tie_guard_I[0].lo ;
 wire \genblk2[0].tie_guard_I[1].lo ;
 wire \genblk2[1].ctrl_ena_buf_I.a ;
 wire \genblk2[1].ctrl_ena_buf_I.z ;
 wire \genblk2[1].pad_ui_in_buf_I[0].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[0].z ;
 wire \genblk2[1].pad_ui_in_buf_I[1].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[1].z ;
 wire \genblk2[1].pad_ui_in_buf_I[2].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[2].z ;
 wire \genblk2[1].pad_ui_in_buf_I[3].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[3].z ;
 wire \genblk2[1].pad_ui_in_buf_I[4].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[4].z ;
 wire \genblk2[1].pad_ui_in_buf_I[5].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[5].z ;
 wire \genblk2[1].pad_ui_in_buf_I[6].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[6].z ;
 wire \genblk2[1].pad_ui_in_buf_I[7].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[7].z ;
 wire \genblk2[1].pad_ui_in_buf_I[8].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[8].z ;
 wire \genblk2[1].pad_ui_in_buf_I[9].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[9].z ;
 wire \genblk2[1].pad_uio_in_buf_I[0].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[0].z ;
 wire \genblk2[1].pad_uio_in_buf_I[1].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[1].z ;
 wire \genblk2[1].pad_uio_in_buf_I[2].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[2].z ;
 wire \genblk2[1].pad_uio_in_buf_I[3].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[3].z ;
 wire \genblk2[1].pad_uio_in_buf_I[4].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[4].z ;
 wire \genblk2[1].pad_uio_in_buf_I[5].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[5].z ;
 wire \genblk2[1].pad_uio_in_buf_I[6].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[6].z ;
 wire \genblk2[1].pad_uio_in_buf_I[7].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[7].z ;
 wire \genblk2[1].sel_cnt_buf_I[0].z ;
 wire \genblk2[1].sel_cnt_buf_I[1].z ;
 wire \genblk2[1].sel_cnt_buf_I[2].z ;
 wire \genblk2[1].sel_cnt_buf_I[3].z ;
 wire \genblk2[1].sel_cnt_buf_I[4].z ;
 wire \genblk2[1].sel_cnt_buf_I[5].z ;
 wire \genblk2[1].sel_cnt_buf_I[6].z ;
 wire \genblk2[1].sel_cnt_buf_I[7].z ;
 wire \genblk2[1].sel_cnt_buf_I[8].z ;
 wire \genblk2[1].tie_guard_I[0].lo ;
 wire \genblk2[1].tie_guard_I[1].lo ;
 wire \sel_cnt_gen[0].cnt_bit_I.d ;
 wire \sel_cnt_gen[1].cnt_bit_I.d ;
 wire \sel_cnt_gen[2].cnt_bit_I.d ;
 wire \sel_cnt_gen[3].cnt_bit_I.d ;
 wire \sel_cnt_gen[4].cnt_bit_I.d ;
 wire \sel_cnt_gen[5].cnt_bit_I.d ;
 wire \sel_cnt_gen[5].cnt_bit_I.q ;
 wire \sel_cnt_gen[6].cnt_bit_I.d ;
 wire \sel_cnt_gen[7].cnt_bit_I.d ;
 wire \sel_cnt_gen[8].cnt_bit_I.d ;
 wire \sel_cnt_gen[9].cnt_bit_I.d ;
 wire \side_ena0_buf_I.a ;
 wire \side_ena0_buf_I.genblk1.l ;
 wire \side_ena1_buf_I.genblk1.l ;
 wire side_sel;
 wire \uio_oe_obuf_I[0].a ;
 wire \uio_oe_obuf_I[0].z ;
 wire \uio_oe_obuf_I[1].a ;
 wire \uio_oe_obuf_I[1].z ;
 wire \uio_oe_obuf_I[2].a ;
 wire \uio_oe_obuf_I[2].z ;
 wire \uio_oe_obuf_I[3].a ;
 wire \uio_oe_obuf_I[3].z ;
 wire \uio_oe_obuf_I[4].a ;
 wire \uio_oe_obuf_I[4].z ;
 wire \uio_oe_obuf_I[5].a ;
 wire \uio_oe_obuf_I[5].z ;
 wire \uio_oe_obuf_I[6].a ;
 wire \uio_oe_obuf_I[6].z ;
 wire \uio_oe_obuf_I[7].a ;
 wire \uio_oe_obuf_I[7].z ;
 wire \uio_oex_ibuf_I[0].z ;
 wire \uio_oex_ibuf_I[10].z ;
 wire \uio_oex_ibuf_I[11].z ;
 wire \uio_oex_ibuf_I[12].z ;
 wire \uio_oex_ibuf_I[13].z ;
 wire \uio_oex_ibuf_I[14].z ;
 wire \uio_oex_ibuf_I[15].z ;
 wire \uio_oex_ibuf_I[1].z ;
 wire \uio_oex_ibuf_I[2].z ;
 wire \uio_oex_ibuf_I[3].z ;
 wire \uio_oex_ibuf_I[4].z ;
 wire \uio_oex_ibuf_I[5].z ;
 wire \uio_oex_ibuf_I[6].z ;
 wire \uio_oex_ibuf_I[7].z ;
 wire \uio_oex_ibuf_I[8].z ;
 wire \uio_oex_ibuf_I[9].z ;
 wire \uio_out_ibuf_I[0].z ;
 wire \uio_out_ibuf_I[10].z ;
 wire \uio_out_ibuf_I[11].z ;
 wire \uio_out_ibuf_I[12].z ;
 wire \uio_out_ibuf_I[13].z ;
 wire \uio_out_ibuf_I[14].z ;
 wire \uio_out_ibuf_I[15].z ;
 wire \uio_out_ibuf_I[1].z ;
 wire \uio_out_ibuf_I[2].z ;
 wire \uio_out_ibuf_I[3].z ;
 wire \uio_out_ibuf_I[4].z ;
 wire \uio_out_ibuf_I[5].z ;
 wire \uio_out_ibuf_I[6].z ;
 wire \uio_out_ibuf_I[7].z ;
 wire \uio_out_ibuf_I[8].z ;
 wire \uio_out_ibuf_I[9].z ;
 wire \uio_out_mux_I[0].x ;
 wire \uio_out_mux_I[1].x ;
 wire \uio_out_mux_I[2].x ;
 wire \uio_out_mux_I[3].x ;
 wire \uio_out_mux_I[4].x ;
 wire \uio_out_mux_I[5].x ;
 wire \uio_out_mux_I[6].x ;
 wire \uio_out_mux_I[7].x ;
 wire \uio_out_obuf_I[0].z ;
 wire \uio_out_obuf_I[1].z ;
 wire \uio_out_obuf_I[2].z ;
 wire \uio_out_obuf_I[3].z ;
 wire \uio_out_obuf_I[4].z ;
 wire \uio_out_obuf_I[5].z ;
 wire \uio_out_obuf_I[6].z ;
 wire \uio_out_obuf_I[7].z ;
 wire \uo_out_ibuf_I[0].z ;
 wire \uo_out_ibuf_I[10].z ;
 wire \uo_out_ibuf_I[11].z ;
 wire \uo_out_ibuf_I[12].z ;
 wire \uo_out_ibuf_I[13].z ;
 wire \uo_out_ibuf_I[14].z ;
 wire \uo_out_ibuf_I[15].z ;
 wire \uo_out_ibuf_I[1].z ;
 wire \uo_out_ibuf_I[2].z ;
 wire \uo_out_ibuf_I[3].z ;
 wire \uo_out_ibuf_I[4].z ;
 wire \uo_out_ibuf_I[5].z ;
 wire \uo_out_ibuf_I[6].z ;
 wire \uo_out_ibuf_I[7].z ;
 wire \uo_out_ibuf_I[8].z ;
 wire \uo_out_ibuf_I[9].z ;
 wire \uo_out_mux_I[0].x ;
 wire \uo_out_mux_I[1].x ;
 wire \uo_out_mux_I[2].x ;
 wire \uo_out_mux_I[3].x ;
 wire \uo_out_mux_I[4].x ;
 wire \uo_out_mux_I[5].x ;
 wire \uo_out_mux_I[6].x ;
 wire \uo_out_mux_I[7].x ;
 wire \uo_out_obuf_I[0].z ;
 wire \uo_out_obuf_I[1].z ;
 wire \uo_out_obuf_I[2].z ;
 wire \uo_out_obuf_I[3].z ;
 wire \uo_out_obuf_I[4].z ;
 wire \uo_out_obuf_I[5].z ;
 wire \uo_out_obuf_I[6].z ;
 wire \uo_out_obuf_I[7].z ;

 sg13g2_inv_1 _0_ (.Y(\genblk1[0].pull ),
    .A(\genblk2[0].ctrl_ena_buf_I.a ));
 sg13g2_inv_1 _1_ (.Y(\genblk1[1].pull ),
    .A(\genblk2[1].ctrl_ena_buf_I.a ));
 sg13g2_antennanp \ctrl_diode_I[0].cell0_I  (.A(ctrl_ena));
 sg13g2_antennanp \ctrl_diode_I[1].cell0_I  (.A(ctrl_sel_inc));
 sg13g2_antennanp \ctrl_diode_I[2].cell0_I  (.A(ctrl_sel_rst_n));
 sg13g2_buf_2 \ctrl_ibuf_I[0].genblk1.cell0_I  (.A(ctrl_ena),
    .X(ctrl_ena_ibuf));
 sg13g2_buf_2 \ctrl_ibuf_I[1].genblk1.cell0_I  (.A(ctrl_sel_inc),
    .X(\ctrl_ibuf_I[1].z ));
 sg13g2_buf_2 \ctrl_ibuf_I[2].genblk1.cell0_I  (.A(ctrl_sel_rst_n),
    .X(\ctrl_ibuf_I[2].z ));
 sg13g2_inv_8 \genblk1[0].tbuf_pol_spine_ow_I.cell0_I  (.Y(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .A(\genblk1[0].pull ));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[1]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[11]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[12]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[13]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[14]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[15]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[16]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[17]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[18]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[19]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[20]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[2]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[21]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[22]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[23]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[24]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[3]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[4]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[5]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[6]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[7]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[8]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[9]));
 sg13g2_ebufn_4 \genblk1[0].tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[10]));
 sg13g2_tielo \genblk1[0].tie_I.genblk1.cell0_I  (.L_LO(\genblk1[0].tbuf_spine_ow_I[0].a ));
 sg13g2_inv_8 \genblk1[1].tbuf_pol_spine_ow_I.cell0_I  (.Y(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .A(\genblk1[1].pull ));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[1]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[11]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[12]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[13]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[14]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[15]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[16]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[17]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[18]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[19]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[20]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[2]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[21]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[22]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[23]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[24]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[3]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[4]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[5]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[6]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[7]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[8]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[9]));
 sg13g2_ebufn_4 \genblk1[1].tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[10]));
 sg13g2_tielo \genblk1[1].tie_I.genblk1.cell0_I  (.L_LO(\genblk1[1].tbuf_spine_ow_I[0].a ));
 sg13g2_buf_8 \genblk2[0].ctrl_ena_buf_I.genblk1.cell0_I  (.A(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].ctrl_ena_buf_I.z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[0].genblk1.cell0_I  (.A(pad_ui_in[0]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[0].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[0].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[0].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[0].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[1].genblk1.cell0_I  (.A(pad_ui_in[1]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[1].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[1].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[1].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[1].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[2].genblk1.cell0_I  (.A(pad_ui_in[2]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[2].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[2].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[2].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[2].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[3].genblk1.cell0_I  (.A(pad_ui_in[3]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[3].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[3].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[3].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[3].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[4].genblk1.cell0_I  (.A(pad_ui_in[4]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[4].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[4].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[4].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[4].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[5].genblk1.cell0_I  (.A(pad_ui_in[5]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[5].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[5].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[5].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[5].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[6].genblk1.cell0_I  (.A(pad_ui_in[6]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[6].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[6].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[6].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[6].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[7].genblk1.cell0_I  (.A(pad_ui_in[7]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[7].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[7].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[7].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[7].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[8].genblk1.cell0_I  (.A(pad_ui_in[8]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[8].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[8].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[8].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[8].z ));
 sg13g2_and2_2 \genblk2[0].pad_ui_in_buf_I[9].genblk1.cell0_I  (.A(pad_ui_in[9]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_ui_in_buf_I[9].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_ui_in_buf_I[9].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[9].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[9].z ));
 sg13g2_and2_2 \genblk2[0].pad_uio_in_buf_I[0].genblk1.cell0_I  (.A(pad_uio_in[0]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_uio_in_buf_I[0].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_uio_in_buf_I[0].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[0].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[0].z ));
 sg13g2_and2_2 \genblk2[0].pad_uio_in_buf_I[1].genblk1.cell0_I  (.A(pad_uio_in[1]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_uio_in_buf_I[1].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_uio_in_buf_I[1].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[1].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[1].z ));
 sg13g2_and2_2 \genblk2[0].pad_uio_in_buf_I[2].genblk1.cell0_I  (.A(pad_uio_in[2]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_uio_in_buf_I[2].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_uio_in_buf_I[2].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[2].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[2].z ));
 sg13g2_and2_2 \genblk2[0].pad_uio_in_buf_I[3].genblk1.cell0_I  (.A(pad_uio_in[3]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_uio_in_buf_I[3].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_uio_in_buf_I[3].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[3].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[3].z ));
 sg13g2_and2_2 \genblk2[0].pad_uio_in_buf_I[4].genblk1.cell0_I  (.A(pad_uio_in[4]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_uio_in_buf_I[4].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_uio_in_buf_I[4].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[4].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[4].z ));
 sg13g2_and2_2 \genblk2[0].pad_uio_in_buf_I[5].genblk1.cell0_I  (.A(pad_uio_in[5]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_uio_in_buf_I[5].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_uio_in_buf_I[5].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[5].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[5].z ));
 sg13g2_and2_2 \genblk2[0].pad_uio_in_buf_I[6].genblk1.cell0_I  (.A(pad_uio_in[6]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_uio_in_buf_I[6].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_uio_in_buf_I[6].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[6].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[6].z ));
 sg13g2_and2_2 \genblk2[0].pad_uio_in_buf_I[7].genblk1.cell0_I  (.A(pad_uio_in[7]),
    .B(\genblk2[0].ctrl_ena_buf_I.a ),
    .X(\genblk2[0].pad_uio_in_buf_I[7].genblk1.l ));
 sg13g2_buf_8 \genblk2[0].pad_uio_in_buf_I[7].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[7].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[7].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[0].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[0].a ),
    .X(\genblk2[0].sel_cnt_buf_I[0].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[1].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[1].a ),
    .X(\genblk2[0].sel_cnt_buf_I[1].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[2].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[2].a ),
    .X(\genblk2[0].sel_cnt_buf_I[2].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[3].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[3].a ),
    .X(\genblk2[0].sel_cnt_buf_I[3].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[4].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[4].a ),
    .X(\genblk2[0].sel_cnt_buf_I[4].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[5].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[5].a ),
    .X(\genblk2[0].sel_cnt_buf_I[5].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[6].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[6].a ),
    .X(\genblk2[0].sel_cnt_buf_I[6].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[7].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[7].a ),
    .X(\genblk2[0].sel_cnt_buf_I[7].z ));
 sg13g2_buf_8 \genblk2[0].sel_cnt_buf_I[8].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[8].a ),
    .X(\genblk2[0].sel_cnt_buf_I[8].z ));
 sg13g2_tielo \genblk2[0].tie_guard_I[0].genblk1.cell0_I  (.L_LO(\genblk2[0].tie_guard_I[0].lo ));
 sg13g2_tielo \genblk2[0].tie_guard_I[1].genblk1.cell0_I  (.L_LO(\genblk2[0].tie_guard_I[1].lo ));
 sg13g2_buf_8 \genblk2[1].ctrl_ena_buf_I.genblk1.cell0_I  (.A(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].ctrl_ena_buf_I.z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[0].genblk1.cell0_I  (.A(pad_ui_in[0]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[0].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[0].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[0].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[0].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[1].genblk1.cell0_I  (.A(pad_ui_in[1]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[1].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[1].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[1].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[1].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[2].genblk1.cell0_I  (.A(pad_ui_in[2]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[2].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[2].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[2].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[2].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[3].genblk1.cell0_I  (.A(pad_ui_in[3]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[3].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[3].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[3].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[3].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[4].genblk1.cell0_I  (.A(pad_ui_in[4]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[4].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[4].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[4].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[4].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[5].genblk1.cell0_I  (.A(pad_ui_in[5]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[5].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[5].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[5].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[5].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[6].genblk1.cell0_I  (.A(pad_ui_in[6]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[6].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[6].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[6].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[6].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[7].genblk1.cell0_I  (.A(pad_ui_in[7]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[7].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[7].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[7].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[7].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[8].genblk1.cell0_I  (.A(pad_ui_in[8]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[8].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[8].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[8].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[8].z ));
 sg13g2_and2_2 \genblk2[1].pad_ui_in_buf_I[9].genblk1.cell0_I  (.A(pad_ui_in[9]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_ui_in_buf_I[9].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_ui_in_buf_I[9].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[9].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[9].z ));
 sg13g2_and2_2 \genblk2[1].pad_uio_in_buf_I[0].genblk1.cell0_I  (.A(pad_uio_in[0]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_uio_in_buf_I[0].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_uio_in_buf_I[0].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[0].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[0].z ));
 sg13g2_and2_2 \genblk2[1].pad_uio_in_buf_I[1].genblk1.cell0_I  (.A(pad_uio_in[1]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_uio_in_buf_I[1].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_uio_in_buf_I[1].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[1].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[1].z ));
 sg13g2_and2_2 \genblk2[1].pad_uio_in_buf_I[2].genblk1.cell0_I  (.A(pad_uio_in[2]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_uio_in_buf_I[2].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_uio_in_buf_I[2].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[2].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[2].z ));
 sg13g2_and2_2 \genblk2[1].pad_uio_in_buf_I[3].genblk1.cell0_I  (.A(pad_uio_in[3]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_uio_in_buf_I[3].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_uio_in_buf_I[3].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[3].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[3].z ));
 sg13g2_and2_2 \genblk2[1].pad_uio_in_buf_I[4].genblk1.cell0_I  (.A(pad_uio_in[4]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_uio_in_buf_I[4].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_uio_in_buf_I[4].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[4].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[4].z ));
 sg13g2_and2_2 \genblk2[1].pad_uio_in_buf_I[5].genblk1.cell0_I  (.A(pad_uio_in[5]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_uio_in_buf_I[5].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_uio_in_buf_I[5].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[5].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[5].z ));
 sg13g2_and2_2 \genblk2[1].pad_uio_in_buf_I[6].genblk1.cell0_I  (.A(pad_uio_in[6]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_uio_in_buf_I[6].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_uio_in_buf_I[6].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[6].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[6].z ));
 sg13g2_and2_2 \genblk2[1].pad_uio_in_buf_I[7].genblk1.cell0_I  (.A(pad_uio_in[7]),
    .B(\genblk2[1].ctrl_ena_buf_I.a ),
    .X(\genblk2[1].pad_uio_in_buf_I[7].genblk1.l ));
 sg13g2_buf_8 \genblk2[1].pad_uio_in_buf_I[7].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[7].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[7].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[0].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[0].a ),
    .X(\genblk2[1].sel_cnt_buf_I[0].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[1].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[1].a ),
    .X(\genblk2[1].sel_cnt_buf_I[1].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[2].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[2].a ),
    .X(\genblk2[1].sel_cnt_buf_I[2].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[3].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[3].a ),
    .X(\genblk2[1].sel_cnt_buf_I[3].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[4].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[4].a ),
    .X(\genblk2[1].sel_cnt_buf_I[4].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[5].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[5].a ),
    .X(\genblk2[1].sel_cnt_buf_I[5].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[6].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[6].a ),
    .X(\genblk2[1].sel_cnt_buf_I[6].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[7].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[7].a ),
    .X(\genblk2[1].sel_cnt_buf_I[7].z ));
 sg13g2_buf_8 \genblk2[1].sel_cnt_buf_I[8].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[8].a ),
    .X(\genblk2[1].sel_cnt_buf_I[8].z ));
 sg13g2_tielo \genblk2[1].tie_guard_I[0].genblk1.cell0_I  (.L_LO(\genblk2[1].tie_guard_I[0].lo ));
 sg13g2_tielo \genblk2[1].tie_guard_I[1].genblk1.cell0_I  (.L_LO(\genblk2[1].tie_guard_I[1].lo ));
 sg13g2_antennanp \pad_ui_in_diode_I[0].cell0_I  (.A(pad_ui_in[0]));
 sg13g2_antennanp \pad_ui_in_diode_I[1].cell0_I  (.A(pad_ui_in[1]));
 sg13g2_antennanp \pad_ui_in_diode_I[2].cell0_I  (.A(pad_ui_in[2]));
 sg13g2_antennanp \pad_ui_in_diode_I[3].cell0_I  (.A(pad_ui_in[3]));
 sg13g2_antennanp \pad_ui_in_diode_I[4].cell0_I  (.A(pad_ui_in[4]));
 sg13g2_antennanp \pad_ui_in_diode_I[5].cell0_I  (.A(pad_ui_in[5]));
 sg13g2_antennanp \pad_ui_in_diode_I[6].cell0_I  (.A(pad_ui_in[6]));
 sg13g2_antennanp \pad_ui_in_diode_I[7].cell0_I  (.A(pad_ui_in[7]));
 sg13g2_antennanp \pad_ui_in_diode_I[8].cell0_I  (.A(pad_ui_in[8]));
 sg13g2_antennanp \pad_ui_in_diode_I[9].cell0_I  (.A(pad_ui_in[9]));
 sg13g2_antennanp \pad_uio_in_diode_I[0].cell0_I  (.A(pad_uio_in[0]));
 sg13g2_antennanp \pad_uio_in_diode_I[1].cell0_I  (.A(pad_uio_in[1]));
 sg13g2_antennanp \pad_uio_in_diode_I[2].cell0_I  (.A(pad_uio_in[2]));
 sg13g2_antennanp \pad_uio_in_diode_I[3].cell0_I  (.A(pad_uio_in[3]));
 sg13g2_antennanp \pad_uio_in_diode_I[4].cell0_I  (.A(pad_uio_in[4]));
 sg13g2_antennanp \pad_uio_in_diode_I[5].cell0_I  (.A(pad_uio_in[5]));
 sg13g2_antennanp \pad_uio_in_diode_I[6].cell0_I  (.A(pad_uio_in[6]));
 sg13g2_antennanp \pad_uio_in_diode_I[7].cell0_I  (.A(pad_uio_in[7]));
 sg13g2_dfrbp_2 \sel_cnt_gen[0].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[0].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[0].a ),
    .Q_N(\sel_cnt_gen[0].cnt_bit_I.d ),
    .CLK(\ctrl_ibuf_I[1].z ));
 sg13g2_dfrbp_2 \sel_cnt_gen[1].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[1].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[1].a ),
    .Q_N(\sel_cnt_gen[1].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[0].cnt_bit_I.d ));
 sg13g2_dfrbp_2 \sel_cnt_gen[2].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[2].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[2].a ),
    .Q_N(\sel_cnt_gen[2].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[1].cnt_bit_I.d ));
 sg13g2_dfrbp_2 \sel_cnt_gen[3].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[3].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[3].a ),
    .Q_N(\sel_cnt_gen[3].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[2].cnt_bit_I.d ));
 sg13g2_dfrbp_2 \sel_cnt_gen[4].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[4].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[4].a ),
    .Q_N(\sel_cnt_gen[4].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[3].cnt_bit_I.d ));
 sg13g2_dfrbp_2 \sel_cnt_gen[5].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[5].cnt_bit_I.d ),
    .Q(\sel_cnt_gen[5].cnt_bit_I.q ),
    .Q_N(\sel_cnt_gen[5].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[4].cnt_bit_I.d ));
 sg13g2_dfrbp_2 \sel_cnt_gen[6].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[6].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[5].a ),
    .Q_N(\sel_cnt_gen[6].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[5].cnt_bit_I.d ));
 sg13g2_dfrbp_2 \sel_cnt_gen[7].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[7].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[6].a ),
    .Q_N(\sel_cnt_gen[7].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[6].cnt_bit_I.d ));
 sg13g2_dfrbp_2 \sel_cnt_gen[8].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[8].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[7].a ),
    .Q_N(\sel_cnt_gen[8].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[7].cnt_bit_I.d ));
 sg13g2_dfrbp_2 \sel_cnt_gen[9].cnt_bit_I.cell0_I  (.RESET_B(\ctrl_ibuf_I[2].z ),
    .D(\sel_cnt_gen[9].cnt_bit_I.d ),
    .Q(\genblk2[0].sel_cnt_buf_I[8].a ),
    .Q_N(\sel_cnt_gen[9].cnt_bit_I.d ),
    .CLK(\sel_cnt_gen[8].cnt_bit_I.d ));
 sg13g2_and2_2 \side_ena0_buf_I.genblk1.cell0_I  (.A(\side_ena0_buf_I.a ),
    .B(ctrl_ena_ibuf),
    .X(\side_ena0_buf_I.genblk1.l ));
 sg13g2_buf_8 \side_ena0_buf_I.genblk1.cell1_I  (.A(\side_ena0_buf_I.genblk1.l ),
    .X(\genblk2[0].ctrl_ena_buf_I.a ));
 sg13g2_inv_2 \side_ena0_gen_I.genblk1.cell0_I  (.Y(\side_ena0_buf_I.a ),
    .A(\sel_cnt_gen[5].cnt_bit_I.q ));
 sg13g2_and2_2 \side_ena1_buf_I.genblk1.cell0_I  (.A(\sel_cnt_gen[5].cnt_bit_I.q ),
    .B(ctrl_ena_ibuf),
    .X(\side_ena1_buf_I.genblk1.l ));
 sg13g2_buf_8 \side_ena1_buf_I.genblk1.cell1_I  (.A(\side_ena1_buf_I.genblk1.l ),
    .X(\genblk2[1].ctrl_ena_buf_I.a ));
 sg13g2_buf_8 \side_sel_buf_I.genblk1.cell0_I  (.A(\sel_cnt_gen[5].cnt_bit_I.q ),
    .X(side_sel));
 sg13g2_antennanp \spine_diode_I[0].cell0_I  (.A(spine_bot_ow[0]));
 sg13g2_antennanp \spine_diode_I[10].cell0_I  (.A(spine_bot_ow[10]));
 sg13g2_antennanp \spine_diode_I[11].cell0_I  (.A(spine_bot_ow[11]));
 sg13g2_antennanp \spine_diode_I[12].cell0_I  (.A(spine_bot_ow[12]));
 sg13g2_antennanp \spine_diode_I[13].cell0_I  (.A(spine_bot_ow[13]));
 sg13g2_antennanp \spine_diode_I[14].cell0_I  (.A(spine_bot_ow[14]));
 sg13g2_antennanp \spine_diode_I[15].cell0_I  (.A(spine_bot_ow[15]));
 sg13g2_antennanp \spine_diode_I[16].cell0_I  (.A(spine_bot_ow[16]));
 sg13g2_antennanp \spine_diode_I[17].cell0_I  (.A(spine_bot_ow[17]));
 sg13g2_antennanp \spine_diode_I[18].cell0_I  (.A(spine_bot_ow[18]));
 sg13g2_antennanp \spine_diode_I[19].cell0_I  (.A(spine_bot_ow[19]));
 sg13g2_antennanp \spine_diode_I[1].cell0_I  (.A(spine_bot_ow[1]));
 sg13g2_antennanp \spine_diode_I[20].cell0_I  (.A(spine_bot_ow[20]));
 sg13g2_antennanp \spine_diode_I[21].cell0_I  (.A(spine_bot_ow[21]));
 sg13g2_antennanp \spine_diode_I[22].cell0_I  (.A(spine_bot_ow[22]));
 sg13g2_antennanp \spine_diode_I[23].cell0_I  (.A(spine_bot_ow[23]));
 sg13g2_antennanp \spine_diode_I[24].cell0_I  (.A(spine_bot_ow[24]));
 sg13g2_antennanp \spine_diode_I[25].cell0_I  (.A(spine_bot_ow[25]));
 sg13g2_antennanp \spine_diode_I[26].cell0_I  (.A(spine_top_ow[0]));
 sg13g2_antennanp \spine_diode_I[27].cell0_I  (.A(spine_top_ow[1]));
 sg13g2_antennanp \spine_diode_I[28].cell0_I  (.A(spine_top_ow[2]));
 sg13g2_antennanp \spine_diode_I[29].cell0_I  (.A(spine_top_ow[3]));
 sg13g2_antennanp \spine_diode_I[2].cell0_I  (.A(spine_bot_ow[2]));
 sg13g2_antennanp \spine_diode_I[30].cell0_I  (.A(spine_top_ow[4]));
 sg13g2_antennanp \spine_diode_I[31].cell0_I  (.A(spine_top_ow[5]));
 sg13g2_antennanp \spine_diode_I[32].cell0_I  (.A(spine_top_ow[6]));
 sg13g2_antennanp \spine_diode_I[33].cell0_I  (.A(spine_top_ow[7]));
 sg13g2_antennanp \spine_diode_I[34].cell0_I  (.A(spine_top_ow[8]));
 sg13g2_antennanp \spine_diode_I[35].cell0_I  (.A(spine_top_ow[9]));
 sg13g2_antennanp \spine_diode_I[36].cell0_I  (.A(spine_top_ow[10]));
 sg13g2_antennanp \spine_diode_I[37].cell0_I  (.A(spine_top_ow[11]));
 sg13g2_antennanp \spine_diode_I[38].cell0_I  (.A(spine_top_ow[12]));
 sg13g2_antennanp \spine_diode_I[39].cell0_I  (.A(spine_top_ow[13]));
 sg13g2_antennanp \spine_diode_I[3].cell0_I  (.A(spine_bot_ow[3]));
 sg13g2_antennanp \spine_diode_I[40].cell0_I  (.A(spine_top_ow[14]));
 sg13g2_antennanp \spine_diode_I[41].cell0_I  (.A(spine_top_ow[15]));
 sg13g2_antennanp \spine_diode_I[42].cell0_I  (.A(spine_top_ow[16]));
 sg13g2_antennanp \spine_diode_I[43].cell0_I  (.A(spine_top_ow[17]));
 sg13g2_antennanp \spine_diode_I[44].cell0_I  (.A(spine_top_ow[18]));
 sg13g2_antennanp \spine_diode_I[45].cell0_I  (.A(spine_top_ow[19]));
 sg13g2_antennanp \spine_diode_I[46].cell0_I  (.A(spine_top_ow[20]));
 sg13g2_antennanp \spine_diode_I[47].cell0_I  (.A(spine_top_ow[21]));
 sg13g2_antennanp \spine_diode_I[48].cell0_I  (.A(spine_top_ow[22]));
 sg13g2_antennanp \spine_diode_I[49].cell0_I  (.A(spine_top_ow[23]));
 sg13g2_antennanp \spine_diode_I[4].cell0_I  (.A(spine_bot_ow[4]));
 sg13g2_antennanp \spine_diode_I[50].cell0_I  (.A(spine_top_ow[24]));
 sg13g2_antennanp \spine_diode_I[51].cell0_I  (.A(spine_top_ow[25]));
 sg13g2_antennanp \spine_diode_I[5].cell0_I  (.A(spine_bot_ow[5]));
 sg13g2_antennanp \spine_diode_I[6].cell0_I  (.A(spine_bot_ow[6]));
 sg13g2_antennanp \spine_diode_I[7].cell0_I  (.A(spine_bot_ow[7]));
 sg13g2_antennanp \spine_diode_I[8].cell0_I  (.A(spine_bot_ow[8]));
 sg13g2_antennanp \spine_diode_I[9].cell0_I  (.A(spine_bot_ow[9]));
 sg13g2_tielo \tie_I.genblk1.cell0_I  (.L_LO(k_zero));
 sg13g2_tiehi \tie_I.genblk2.cell1_I  (.L_HI(k_one));
 sg13g2_inv_8 \uio_oe_obuf_I[0].genblk1.cell0_I  (.Y(\uio_oe_obuf_I[0].z ),
    .A(\uio_oe_obuf_I[0].a ));
 sg13g2_inv_8 \uio_oe_obuf_I[1].genblk1.cell0_I  (.Y(\uio_oe_obuf_I[1].z ),
    .A(\uio_oe_obuf_I[1].a ));
 sg13g2_inv_8 \uio_oe_obuf_I[2].genblk1.cell0_I  (.Y(\uio_oe_obuf_I[2].z ),
    .A(\uio_oe_obuf_I[2].a ));
 sg13g2_inv_8 \uio_oe_obuf_I[3].genblk1.cell0_I  (.Y(\uio_oe_obuf_I[3].z ),
    .A(\uio_oe_obuf_I[3].a ));
 sg13g2_inv_8 \uio_oe_obuf_I[4].genblk1.cell0_I  (.Y(\uio_oe_obuf_I[4].z ),
    .A(\uio_oe_obuf_I[4].a ));
 sg13g2_inv_8 \uio_oe_obuf_I[5].genblk1.cell0_I  (.Y(\uio_oe_obuf_I[5].z ),
    .A(\uio_oe_obuf_I[5].a ));
 sg13g2_inv_8 \uio_oe_obuf_I[6].genblk1.cell0_I  (.Y(\uio_oe_obuf_I[6].z ),
    .A(\uio_oe_obuf_I[6].a ));
 sg13g2_inv_8 \uio_oe_obuf_I[7].genblk1.cell0_I  (.Y(\uio_oe_obuf_I[7].z ),
    .A(\uio_oe_obuf_I[7].a ));
 sg13g2_inv_2 \uio_oex_ibuf_I[0].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[0].z ),
    .A(spine_bot_ow[17]));
 sg13g2_inv_2 \uio_oex_ibuf_I[10].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[10].z ),
    .A(spine_top_ow[19]));
 sg13g2_inv_2 \uio_oex_ibuf_I[11].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[11].z ),
    .A(spine_top_ow[20]));
 sg13g2_inv_2 \uio_oex_ibuf_I[12].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[12].z ),
    .A(spine_top_ow[21]));
 sg13g2_inv_2 \uio_oex_ibuf_I[13].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[13].z ),
    .A(spine_top_ow[22]));
 sg13g2_inv_2 \uio_oex_ibuf_I[14].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[14].z ),
    .A(spine_top_ow[23]));
 sg13g2_inv_2 \uio_oex_ibuf_I[15].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[15].z ),
    .A(spine_top_ow[24]));
 sg13g2_inv_2 \uio_oex_ibuf_I[1].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[1].z ),
    .A(spine_bot_ow[18]));
 sg13g2_inv_2 \uio_oex_ibuf_I[2].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[2].z ),
    .A(spine_bot_ow[19]));
 sg13g2_inv_2 \uio_oex_ibuf_I[3].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[3].z ),
    .A(spine_bot_ow[20]));
 sg13g2_inv_2 \uio_oex_ibuf_I[4].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[4].z ),
    .A(spine_bot_ow[21]));
 sg13g2_inv_2 \uio_oex_ibuf_I[5].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[5].z ),
    .A(spine_bot_ow[22]));
 sg13g2_inv_2 \uio_oex_ibuf_I[6].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[6].z ),
    .A(spine_bot_ow[23]));
 sg13g2_inv_2 \uio_oex_ibuf_I[7].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[7].z ),
    .A(spine_bot_ow[24]));
 sg13g2_inv_2 \uio_oex_ibuf_I[8].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[8].z ),
    .A(spine_top_ow[17]));
 sg13g2_inv_2 \uio_oex_ibuf_I[9].genblk1.cell0_I  (.Y(\uio_oex_ibuf_I[9].z ),
    .A(spine_top_ow[18]));
 sg13g2_mux2_1 \uio_oex_mux_I[0].cell0_I  (.A0(\uio_oex_ibuf_I[0].z ),
    .A1(\uio_oex_ibuf_I[8].z ),
    .S(side_sel),
    .X(\uio_oe_obuf_I[0].a ));
 sg13g2_mux2_1 \uio_oex_mux_I[1].cell0_I  (.A0(\uio_oex_ibuf_I[1].z ),
    .A1(\uio_oex_ibuf_I[9].z ),
    .S(side_sel),
    .X(\uio_oe_obuf_I[1].a ));
 sg13g2_mux2_1 \uio_oex_mux_I[2].cell0_I  (.A0(\uio_oex_ibuf_I[2].z ),
    .A1(\uio_oex_ibuf_I[10].z ),
    .S(side_sel),
    .X(\uio_oe_obuf_I[2].a ));
 sg13g2_mux2_1 \uio_oex_mux_I[3].cell0_I  (.A0(\uio_oex_ibuf_I[3].z ),
    .A1(\uio_oex_ibuf_I[11].z ),
    .S(side_sel),
    .X(\uio_oe_obuf_I[3].a ));
 sg13g2_mux2_1 \uio_oex_mux_I[4].cell0_I  (.A0(\uio_oex_ibuf_I[4].z ),
    .A1(\uio_oex_ibuf_I[12].z ),
    .S(side_sel),
    .X(\uio_oe_obuf_I[4].a ));
 sg13g2_mux2_1 \uio_oex_mux_I[5].cell0_I  (.A0(\uio_oex_ibuf_I[5].z ),
    .A1(\uio_oex_ibuf_I[13].z ),
    .S(side_sel),
    .X(\uio_oe_obuf_I[5].a ));
 sg13g2_mux2_1 \uio_oex_mux_I[6].cell0_I  (.A0(\uio_oex_ibuf_I[6].z ),
    .A1(\uio_oex_ibuf_I[14].z ),
    .S(side_sel),
    .X(\uio_oe_obuf_I[6].a ));
 sg13g2_mux2_1 \uio_oex_mux_I[7].cell0_I  (.A0(\uio_oex_ibuf_I[7].z ),
    .A1(\uio_oex_ibuf_I[15].z ),
    .S(side_sel),
    .X(\uio_oe_obuf_I[7].a ));
 sg13g2_inv_2 \uio_out_ibuf_I[0].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[0].z ),
    .A(spine_bot_ow[9]));
 sg13g2_inv_2 \uio_out_ibuf_I[10].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[10].z ),
    .A(spine_top_ow[11]));
 sg13g2_inv_2 \uio_out_ibuf_I[11].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[11].z ),
    .A(spine_top_ow[12]));
 sg13g2_inv_2 \uio_out_ibuf_I[12].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[12].z ),
    .A(spine_top_ow[13]));
 sg13g2_inv_2 \uio_out_ibuf_I[13].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[13].z ),
    .A(spine_top_ow[14]));
 sg13g2_inv_2 \uio_out_ibuf_I[14].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[14].z ),
    .A(spine_top_ow[15]));
 sg13g2_inv_2 \uio_out_ibuf_I[15].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[15].z ),
    .A(spine_top_ow[16]));
 sg13g2_inv_2 \uio_out_ibuf_I[1].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[1].z ),
    .A(spine_bot_ow[10]));
 sg13g2_inv_2 \uio_out_ibuf_I[2].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[2].z ),
    .A(spine_bot_ow[11]));
 sg13g2_inv_2 \uio_out_ibuf_I[3].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[3].z ),
    .A(spine_bot_ow[12]));
 sg13g2_inv_2 \uio_out_ibuf_I[4].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[4].z ),
    .A(spine_bot_ow[13]));
 sg13g2_inv_2 \uio_out_ibuf_I[5].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[5].z ),
    .A(spine_bot_ow[14]));
 sg13g2_inv_2 \uio_out_ibuf_I[6].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[6].z ),
    .A(spine_bot_ow[15]));
 sg13g2_inv_2 \uio_out_ibuf_I[7].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[7].z ),
    .A(spine_bot_ow[16]));
 sg13g2_inv_2 \uio_out_ibuf_I[8].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[8].z ),
    .A(spine_top_ow[9]));
 sg13g2_inv_2 \uio_out_ibuf_I[9].genblk1.cell0_I  (.Y(\uio_out_ibuf_I[9].z ),
    .A(spine_top_ow[10]));
 sg13g2_mux2_1 \uio_out_mux_I[0].cell0_I  (.A0(\uio_out_ibuf_I[0].z ),
    .A1(\uio_out_ibuf_I[8].z ),
    .S(side_sel),
    .X(\uio_out_mux_I[0].x ));
 sg13g2_mux2_1 \uio_out_mux_I[1].cell0_I  (.A0(\uio_out_ibuf_I[1].z ),
    .A1(\uio_out_ibuf_I[9].z ),
    .S(side_sel),
    .X(\uio_out_mux_I[1].x ));
 sg13g2_mux2_1 \uio_out_mux_I[2].cell0_I  (.A0(\uio_out_ibuf_I[2].z ),
    .A1(\uio_out_ibuf_I[10].z ),
    .S(side_sel),
    .X(\uio_out_mux_I[2].x ));
 sg13g2_mux2_1 \uio_out_mux_I[3].cell0_I  (.A0(\uio_out_ibuf_I[3].z ),
    .A1(\uio_out_ibuf_I[11].z ),
    .S(side_sel),
    .X(\uio_out_mux_I[3].x ));
 sg13g2_mux2_1 \uio_out_mux_I[4].cell0_I  (.A0(\uio_out_ibuf_I[4].z ),
    .A1(\uio_out_ibuf_I[12].z ),
    .S(side_sel),
    .X(\uio_out_mux_I[4].x ));
 sg13g2_mux2_1 \uio_out_mux_I[5].cell0_I  (.A0(\uio_out_ibuf_I[5].z ),
    .A1(\uio_out_ibuf_I[13].z ),
    .S(side_sel),
    .X(\uio_out_mux_I[5].x ));
 sg13g2_mux2_1 \uio_out_mux_I[6].cell0_I  (.A0(\uio_out_ibuf_I[6].z ),
    .A1(\uio_out_ibuf_I[14].z ),
    .S(side_sel),
    .X(\uio_out_mux_I[6].x ));
 sg13g2_mux2_1 \uio_out_mux_I[7].cell0_I  (.A0(\uio_out_ibuf_I[7].z ),
    .A1(\uio_out_ibuf_I[15].z ),
    .S(side_sel),
    .X(\uio_out_mux_I[7].x ));
 sg13g2_inv_8 \uio_out_obuf_I[0].genblk1.cell0_I  (.Y(\uio_out_obuf_I[0].z ),
    .A(\uio_out_mux_I[0].x ));
 sg13g2_inv_8 \uio_out_obuf_I[1].genblk1.cell0_I  (.Y(\uio_out_obuf_I[1].z ),
    .A(\uio_out_mux_I[1].x ));
 sg13g2_inv_8 \uio_out_obuf_I[2].genblk1.cell0_I  (.Y(\uio_out_obuf_I[2].z ),
    .A(\uio_out_mux_I[2].x ));
 sg13g2_inv_8 \uio_out_obuf_I[3].genblk1.cell0_I  (.Y(\uio_out_obuf_I[3].z ),
    .A(\uio_out_mux_I[3].x ));
 sg13g2_inv_8 \uio_out_obuf_I[4].genblk1.cell0_I  (.Y(\uio_out_obuf_I[4].z ),
    .A(\uio_out_mux_I[4].x ));
 sg13g2_inv_8 \uio_out_obuf_I[5].genblk1.cell0_I  (.Y(\uio_out_obuf_I[5].z ),
    .A(\uio_out_mux_I[5].x ));
 sg13g2_inv_8 \uio_out_obuf_I[6].genblk1.cell0_I  (.Y(\uio_out_obuf_I[6].z ),
    .A(\uio_out_mux_I[6].x ));
 sg13g2_inv_8 \uio_out_obuf_I[7].genblk1.cell0_I  (.Y(\uio_out_obuf_I[7].z ),
    .A(\uio_out_mux_I[7].x ));
 sg13g2_inv_2 \uo_out_ibuf_I[0].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[0].z ),
    .A(spine_bot_ow[1]));
 sg13g2_inv_2 \uo_out_ibuf_I[10].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[10].z ),
    .A(spine_top_ow[3]));
 sg13g2_inv_2 \uo_out_ibuf_I[11].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[11].z ),
    .A(spine_top_ow[4]));
 sg13g2_inv_2 \uo_out_ibuf_I[12].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[12].z ),
    .A(spine_top_ow[5]));
 sg13g2_inv_2 \uo_out_ibuf_I[13].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[13].z ),
    .A(spine_top_ow[6]));
 sg13g2_inv_2 \uo_out_ibuf_I[14].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[14].z ),
    .A(spine_top_ow[7]));
 sg13g2_inv_2 \uo_out_ibuf_I[15].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[15].z ),
    .A(spine_top_ow[8]));
 sg13g2_inv_2 \uo_out_ibuf_I[1].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[1].z ),
    .A(spine_bot_ow[2]));
 sg13g2_inv_2 \uo_out_ibuf_I[2].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[2].z ),
    .A(spine_bot_ow[3]));
 sg13g2_inv_2 \uo_out_ibuf_I[3].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[3].z ),
    .A(spine_bot_ow[4]));
 sg13g2_inv_2 \uo_out_ibuf_I[4].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[4].z ),
    .A(spine_bot_ow[5]));
 sg13g2_inv_2 \uo_out_ibuf_I[5].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[5].z ),
    .A(spine_bot_ow[6]));
 sg13g2_inv_2 \uo_out_ibuf_I[6].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[6].z ),
    .A(spine_bot_ow[7]));
 sg13g2_inv_2 \uo_out_ibuf_I[7].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[7].z ),
    .A(spine_bot_ow[8]));
 sg13g2_inv_2 \uo_out_ibuf_I[8].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[8].z ),
    .A(spine_top_ow[1]));
 sg13g2_inv_2 \uo_out_ibuf_I[9].genblk1.cell0_I  (.Y(\uo_out_ibuf_I[9].z ),
    .A(spine_top_ow[2]));
 sg13g2_mux2_1 \uo_out_mux_I[0].cell0_I  (.A0(\uo_out_ibuf_I[0].z ),
    .A1(\uo_out_ibuf_I[8].z ),
    .S(side_sel),
    .X(\uo_out_mux_I[0].x ));
 sg13g2_mux2_1 \uo_out_mux_I[1].cell0_I  (.A0(\uo_out_ibuf_I[1].z ),
    .A1(\uo_out_ibuf_I[9].z ),
    .S(side_sel),
    .X(\uo_out_mux_I[1].x ));
 sg13g2_mux2_1 \uo_out_mux_I[2].cell0_I  (.A0(\uo_out_ibuf_I[2].z ),
    .A1(\uo_out_ibuf_I[10].z ),
    .S(side_sel),
    .X(\uo_out_mux_I[2].x ));
 sg13g2_mux2_1 \uo_out_mux_I[3].cell0_I  (.A0(\uo_out_ibuf_I[3].z ),
    .A1(\uo_out_ibuf_I[11].z ),
    .S(side_sel),
    .X(\uo_out_mux_I[3].x ));
 sg13g2_mux2_1 \uo_out_mux_I[4].cell0_I  (.A0(\uo_out_ibuf_I[4].z ),
    .A1(\uo_out_ibuf_I[12].z ),
    .S(side_sel),
    .X(\uo_out_mux_I[4].x ));
 sg13g2_mux2_1 \uo_out_mux_I[5].cell0_I  (.A0(\uo_out_ibuf_I[5].z ),
    .A1(\uo_out_ibuf_I[13].z ),
    .S(side_sel),
    .X(\uo_out_mux_I[5].x ));
 sg13g2_mux2_1 \uo_out_mux_I[6].cell0_I  (.A0(\uo_out_ibuf_I[6].z ),
    .A1(\uo_out_ibuf_I[14].z ),
    .S(side_sel),
    .X(\uo_out_mux_I[6].x ));
 sg13g2_mux2_1 \uo_out_mux_I[7].cell0_I  (.A0(\uo_out_ibuf_I[7].z ),
    .A1(\uo_out_ibuf_I[15].z ),
    .S(side_sel),
    .X(\uo_out_mux_I[7].x ));
 sg13g2_inv_8 \uo_out_obuf_I[0].genblk1.cell0_I  (.Y(\uo_out_obuf_I[0].z ),
    .A(\uo_out_mux_I[0].x ));
 sg13g2_inv_8 \uo_out_obuf_I[1].genblk1.cell0_I  (.Y(\uo_out_obuf_I[1].z ),
    .A(\uo_out_mux_I[1].x ));
 sg13g2_inv_8 \uo_out_obuf_I[2].genblk1.cell0_I  (.Y(\uo_out_obuf_I[2].z ),
    .A(\uo_out_mux_I[2].x ));
 sg13g2_inv_8 \uo_out_obuf_I[3].genblk1.cell0_I  (.Y(\uo_out_obuf_I[3].z ),
    .A(\uo_out_mux_I[3].x ));
 sg13g2_inv_8 \uo_out_obuf_I[4].genblk1.cell0_I  (.Y(\uo_out_obuf_I[4].z ),
    .A(\uo_out_mux_I[4].x ));
 sg13g2_inv_8 \uo_out_obuf_I[5].genblk1.cell0_I  (.Y(\uo_out_obuf_I[5].z ),
    .A(\uo_out_mux_I[5].x ));
 sg13g2_inv_8 \uo_out_obuf_I[6].genblk1.cell0_I  (.Y(\uo_out_obuf_I[6].z ),
    .A(\uo_out_mux_I[6].x ));
 sg13g2_inv_8 \uo_out_obuf_I[7].genblk1.cell0_I  (.Y(\uo_out_obuf_I[7].z ),
    .A(\uo_out_mux_I[7].x ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_4 FILLER_0_28 ();
 sg13g2_fill_1 FILLER_0_32 ();
 sg13g2_decap_8 FILLER_0_36 ();
 sg13g2_decap_8 FILLER_0_43 ();
 sg13g2_decap_8 FILLER_0_50 ();
 sg13g2_decap_4 FILLER_0_57 ();
 sg13g2_fill_1 FILLER_0_61 ();
 sg13g2_fill_2 FILLER_0_65 ();
 sg13g2_decap_4 FILLER_0_70 ();
 sg13g2_fill_2 FILLER_0_74 ();
 sg13g2_fill_1 FILLER_0_79 ();
 sg13g2_decap_8 FILLER_0_83 ();
 sg13g2_decap_8 FILLER_0_90 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_4 FILLER_0_117 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_141 ();
 sg13g2_decap_8 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_155 ();
 sg13g2_fill_1 FILLER_0_162 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_8 FILLER_0_180 ();
 sg13g2_fill_1 FILLER_0_187 ();
 sg13g2_decap_4 FILLER_1_0 ();
 sg13g2_decap_4 FILLER_1_46 ();
 sg13g2_fill_1 FILLER_1_50 ();
 sg13g2_fill_2 FILLER_1_66 ();
 sg13g2_fill_1 FILLER_1_81 ();
 sg13g2_fill_1 FILLER_1_91 ();
 sg13g2_fill_2 FILLER_1_96 ();
 sg13g2_fill_1 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_132 ();
 sg13g2_fill_2 FILLER_1_139 ();
 sg13g2_fill_1 FILLER_1_141 ();
 sg13g2_fill_2 FILLER_1_159 ();
 sg13g2_fill_1 FILLER_1_161 ();
 sg13g2_decap_4 FILLER_1_182 ();
 sg13g2_fill_2 FILLER_1_186 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_1 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_32 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_fill_1 FILLER_2_92 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_4 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_122 ();
 sg13g2_fill_2 FILLER_2_135 ();
 sg13g2_fill_1 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_fill_2 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_10 ();
 sg13g2_decap_8 FILLER_3_17 ();
 sg13g2_decap_4 FILLER_3_24 ();
 sg13g2_decap_8 FILLER_3_36 ();
 sg13g2_decap_4 FILLER_3_43 ();
 sg13g2_fill_1 FILLER_3_47 ();
 sg13g2_decap_4 FILLER_3_63 ();
 sg13g2_fill_2 FILLER_3_67 ();
 sg13g2_decap_4 FILLER_3_73 ();
 sg13g2_fill_1 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_82 ();
 sg13g2_decap_8 FILLER_3_89 ();
 sg13g2_decap_8 FILLER_3_96 ();
 sg13g2_decap_8 FILLER_3_103 ();
 sg13g2_decap_8 FILLER_3_110 ();
 sg13g2_decap_8 FILLER_3_117 ();
 sg13g2_decap_8 FILLER_3_124 ();
 sg13g2_decap_8 FILLER_3_131 ();
 sg13g2_decap_8 FILLER_3_166 ();
 sg13g2_decap_8 FILLER_3_173 ();
 sg13g2_decap_8 FILLER_3_180 ();
 sg13g2_fill_1 FILLER_3_187 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_30 ();
 sg13g2_decap_8 FILLER_4_34 ();
 sg13g2_decap_8 FILLER_4_41 ();
 sg13g2_decap_8 FILLER_4_48 ();
 sg13g2_decap_8 FILLER_4_55 ();
 sg13g2_fill_2 FILLER_4_62 ();
 sg13g2_fill_1 FILLER_4_64 ();
 sg13g2_decap_4 FILLER_4_80 ();
 sg13g2_fill_2 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_100 ();
 sg13g2_fill_1 FILLER_4_107 ();
 sg13g2_decap_4 FILLER_4_134 ();
 sg13g2_fill_2 FILLER_4_138 ();
 sg13g2_decap_8 FILLER_4_146 ();
 sg13g2_decap_4 FILLER_4_153 ();
 sg13g2_decap_4 FILLER_4_167 ();
 sg13g2_fill_1 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_4 FILLER_4_182 ();
 sg13g2_fill_2 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_10 ();
 sg13g2_decap_8 FILLER_5_17 ();
 sg13g2_fill_2 FILLER_5_24 ();
 sg13g2_decap_8 FILLER_5_41 ();
 sg13g2_decap_8 FILLER_5_48 ();
 sg13g2_decap_8 FILLER_5_55 ();
 sg13g2_decap_8 FILLER_5_62 ();
 sg13g2_decap_8 FILLER_5_69 ();
 sg13g2_decap_8 FILLER_5_76 ();
 sg13g2_decap_8 FILLER_5_83 ();
 sg13g2_decap_8 FILLER_5_90 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_fill_1 FILLER_5_104 ();
 sg13g2_decap_8 FILLER_5_124 ();
 sg13g2_decap_8 FILLER_5_131 ();
 sg13g2_decap_4 FILLER_5_138 ();
 sg13g2_decap_8 FILLER_5_155 ();
 sg13g2_decap_8 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_169 ();
 sg13g2_fill_2 FILLER_5_176 ();
 sg13g2_decap_8 FILLER_5_181 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_fill_2 FILLER_6_35 ();
 sg13g2_fill_1 FILLER_6_37 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_60 ();
 sg13g2_decap_4 FILLER_6_76 ();
 sg13g2_fill_1 FILLER_6_80 ();
 sg13g2_decap_8 FILLER_6_85 ();
 sg13g2_fill_2 FILLER_6_97 ();
 sg13g2_fill_1 FILLER_6_99 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_fill_2 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_150 ();
 sg13g2_decap_4 FILLER_6_157 ();
 sg13g2_decap_8 FILLER_6_171 ();
 sg13g2_decap_8 FILLER_6_178 ();
 sg13g2_fill_2 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_187 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_11 ();
 sg13g2_fill_1 FILLER_7_18 ();
 sg13g2_fill_1 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_53 ();
 sg13g2_decap_4 FILLER_7_60 ();
 sg13g2_decap_4 FILLER_7_79 ();
 sg13g2_fill_1 FILLER_7_83 ();
 sg13g2_decap_8 FILLER_7_94 ();
 sg13g2_decap_8 FILLER_7_101 ();
 sg13g2_decap_8 FILLER_7_108 ();
 sg13g2_decap_8 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_152 ();
 sg13g2_fill_1 FILLER_7_159 ();
 sg13g2_decap_8 FILLER_7_170 ();
 sg13g2_decap_8 FILLER_7_177 ();
 sg13g2_decap_4 FILLER_7_184 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_fill_1 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_26 ();
 sg13g2_decap_8 FILLER_8_33 ();
 sg13g2_decap_8 FILLER_8_40 ();
 sg13g2_fill_1 FILLER_8_47 ();
 sg13g2_fill_2 FILLER_8_63 ();
 sg13g2_fill_2 FILLER_8_80 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_decap_8 FILLER_8_97 ();
 sg13g2_decap_8 FILLER_8_104 ();
 sg13g2_decap_8 FILLER_8_111 ();
 sg13g2_decap_8 FILLER_8_118 ();
 sg13g2_decap_8 FILLER_8_125 ();
 sg13g2_decap_4 FILLER_8_132 ();
 sg13g2_decap_4 FILLER_8_155 ();
 sg13g2_decap_8 FILLER_8_169 ();
 sg13g2_decap_8 FILLER_8_176 ();
 sg13g2_decap_4 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_36 ();
 sg13g2_decap_4 FILLER_9_43 ();
 sg13g2_decap_8 FILLER_9_62 ();
 sg13g2_decap_8 FILLER_9_69 ();
 sg13g2_decap_8 FILLER_9_76 ();
 sg13g2_fill_1 FILLER_9_87 ();
 sg13g2_decap_4 FILLER_9_98 ();
 sg13g2_fill_2 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_169 ();
 sg13g2_decap_8 FILLER_9_176 ();
 sg13g2_decap_4 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_187 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_77 ();
 sg13g2_fill_1 FILLER_10_79 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_4 FILLER_10_95 ();
 sg13g2_fill_1 FILLER_10_99 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_4 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_157 ();
 sg13g2_decap_8 FILLER_10_164 ();
 sg13g2_decap_8 FILLER_10_171 ();
 sg13g2_decap_8 FILLER_10_178 ();
 sg13g2_fill_2 FILLER_10_185 ();
 sg13g2_fill_1 FILLER_10_187 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_44 ();
 sg13g2_fill_2 FILLER_11_51 ();
 sg13g2_decap_8 FILLER_11_68 ();
 sg13g2_fill_2 FILLER_11_75 ();
 sg13g2_fill_1 FILLER_11_80 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_91 ();
 sg13g2_fill_1 FILLER_11_93 ();
 sg13g2_decap_8 FILLER_11_106 ();
 sg13g2_decap_8 FILLER_11_113 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_decap_8 FILLER_11_157 ();
 sg13g2_decap_8 FILLER_11_164 ();
 sg13g2_decap_8 FILLER_11_171 ();
 sg13g2_decap_8 FILLER_11_178 ();
 sg13g2_fill_2 FILLER_11_185 ();
 sg13g2_fill_1 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_11 ();
 sg13g2_fill_2 FILLER_12_15 ();
 sg13g2_fill_2 FILLER_12_20 ();
 sg13g2_decap_4 FILLER_12_52 ();
 sg13g2_fill_2 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_73 ();
 sg13g2_decap_4 FILLER_12_80 ();
 sg13g2_decap_8 FILLER_12_97 ();
 sg13g2_decap_8 FILLER_12_104 ();
 sg13g2_decap_8 FILLER_12_111 ();
 sg13g2_decap_8 FILLER_12_118 ();
 sg13g2_decap_8 FILLER_12_125 ();
 sg13g2_decap_8 FILLER_12_132 ();
 sg13g2_decap_4 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_fill_2 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_4 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_18 ();
 sg13g2_decap_4 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_39 ();
 sg13g2_fill_2 FILLER_13_55 ();
 sg13g2_fill_1 FILLER_13_57 ();
 sg13g2_decap_8 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_106 ();
 sg13g2_fill_1 FILLER_13_108 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_fill_2 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_fill_2 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_decap_8 FILLER_14_86 ();
 sg13g2_decap_8 FILLER_14_93 ();
 sg13g2_decap_8 FILLER_14_100 ();
 sg13g2_fill_2 FILLER_14_107 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_fill_1 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_fill_2 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_22 ();
 sg13g2_decap_4 FILLER_15_29 ();
 sg13g2_fill_2 FILLER_15_33 ();
 sg13g2_decap_8 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_48 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_fill_2 FILLER_15_67 ();
 sg13g2_fill_1 FILLER_15_69 ();
 sg13g2_fill_2 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_76 ();
 sg13g2_decap_8 FILLER_15_87 ();
 sg13g2_fill_2 FILLER_15_94 ();
 sg13g2_decap_8 FILLER_15_121 ();
 sg13g2_decap_8 FILLER_15_128 ();
 sg13g2_decap_8 FILLER_15_135 ();
 sg13g2_decap_8 FILLER_15_142 ();
 sg13g2_decap_8 FILLER_15_149 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_decap_8 FILLER_15_163 ();
 sg13g2_decap_8 FILLER_15_170 ();
 sg13g2_decap_8 FILLER_15_177 ();
 sg13g2_decap_4 FILLER_15_184 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_19 ();
 sg13g2_fill_2 FILLER_16_30 ();
 sg13g2_fill_2 FILLER_16_38 ();
 sg13g2_fill_1 FILLER_16_43 ();
 sg13g2_fill_1 FILLER_16_48 ();
 sg13g2_fill_1 FILLER_16_52 ();
 sg13g2_fill_2 FILLER_16_57 ();
 sg13g2_fill_1 FILLER_16_59 ();
 sg13g2_fill_2 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_65 ();
 sg13g2_decap_4 FILLER_16_69 ();
 sg13g2_decap_8 FILLER_16_76 ();
 sg13g2_decap_8 FILLER_16_83 ();
 sg13g2_fill_2 FILLER_16_90 ();
 sg13g2_fill_1 FILLER_16_92 ();
 sg13g2_decap_8 FILLER_16_106 ();
 sg13g2_decap_8 FILLER_16_113 ();
 sg13g2_decap_8 FILLER_16_120 ();
 sg13g2_decap_8 FILLER_16_127 ();
 sg13g2_decap_8 FILLER_16_134 ();
 sg13g2_decap_4 FILLER_16_141 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_18 ();
 sg13g2_fill_1 FILLER_17_24 ();
 sg13g2_decap_8 FILLER_17_32 ();
 sg13g2_fill_2 FILLER_17_39 ();
 sg13g2_fill_2 FILLER_17_51 ();
 sg13g2_fill_1 FILLER_17_53 ();
 sg13g2_decap_8 FILLER_17_62 ();
 sg13g2_decap_8 FILLER_17_69 ();
 sg13g2_decap_8 FILLER_17_76 ();
 sg13g2_fill_2 FILLER_17_83 ();
 sg13g2_decap_8 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_decap_4 FILLER_17_116 ();
 sg13g2_decap_8 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_4 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_27 ();
 sg13g2_decap_8 FILLER_18_34 ();
 sg13g2_decap_8 FILLER_18_41 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_67 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_4 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_4 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_45 ();
 sg13g2_decap_8 FILLER_19_125 ();
 sg13g2_decap_8 FILLER_19_132 ();
 sg13g2_decap_8 FILLER_19_139 ();
 sg13g2_decap_8 FILLER_19_146 ();
 sg13g2_decap_8 FILLER_19_153 ();
 sg13g2_decap_8 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_4 FILLER_20_53 ();
 sg13g2_fill_1 FILLER_20_57 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_fill_2 FILLER_20_130 ();
 sg13g2_fill_1 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_146 ();
 sg13g2_decap_8 FILLER_20_153 ();
 sg13g2_decap_8 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_decap_8 FILLER_20_174 ();
 sg13g2_decap_8 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_fill_2 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_52 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_decap_4 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_decap_8 FILLER_21_96 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_44 ();
 sg13g2_decap_8 FILLER_22_51 ();
 sg13g2_decap_8 FILLER_22_58 ();
 sg13g2_decap_8 FILLER_22_65 ();
 sg13g2_decap_8 FILLER_22_72 ();
 sg13g2_decap_8 FILLER_22_79 ();
 sg13g2_decap_8 FILLER_22_86 ();
 sg13g2_decap_8 FILLER_22_93 ();
 sg13g2_decap_8 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_107 ();
 sg13g2_decap_8 FILLER_22_114 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_decap_8 FILLER_22_128 ();
 sg13g2_decap_4 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_152 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_187 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_36 ();
 sg13g2_fill_2 FILLER_23_40 ();
 sg13g2_decap_8 FILLER_23_52 ();
 sg13g2_decap_8 FILLER_23_59 ();
 sg13g2_decap_8 FILLER_23_66 ();
 sg13g2_decap_8 FILLER_23_73 ();
 sg13g2_decap_8 FILLER_23_80 ();
 sg13g2_decap_8 FILLER_23_87 ();
 sg13g2_decap_8 FILLER_23_94 ();
 sg13g2_decap_8 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_115 ();
 sg13g2_decap_8 FILLER_23_122 ();
 sg13g2_decap_8 FILLER_23_129 ();
 sg13g2_decap_8 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_156 ();
 sg13g2_decap_8 FILLER_23_163 ();
 sg13g2_decap_8 FILLER_23_170 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_decap_4 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_25 ();
 sg13g2_decap_4 FILLER_24_55 ();
 sg13g2_fill_1 FILLER_24_59 ();
 sg13g2_fill_2 FILLER_24_63 ();
 sg13g2_decap_4 FILLER_24_68 ();
 sg13g2_fill_2 FILLER_24_72 ();
 sg13g2_decap_8 FILLER_24_89 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_decap_4 FILLER_24_103 ();
 sg13g2_fill_1 FILLER_24_107 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_fill_2 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_187 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_47 ();
 sg13g2_decap_8 FILLER_25_54 ();
 sg13g2_decap_4 FILLER_25_61 ();
 sg13g2_fill_1 FILLER_25_65 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_75 ();
 sg13g2_decap_4 FILLER_25_82 ();
 sg13g2_fill_1 FILLER_25_86 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_46 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_2 FILLER_26_93 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_4 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_83 ();
 sg13g2_decap_8 FILLER_27_90 ();
 sg13g2_decap_8 FILLER_27_97 ();
 sg13g2_decap_8 FILLER_27_104 ();
 sg13g2_decap_8 FILLER_27_111 ();
 sg13g2_decap_8 FILLER_27_118 ();
 sg13g2_decap_8 FILLER_27_125 ();
 sg13g2_fill_2 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_134 ();
 sg13g2_decap_8 FILLER_27_148 ();
 sg13g2_decap_4 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_170 ();
 sg13g2_decap_8 FILLER_27_177 ();
 sg13g2_decap_4 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_33 ();
 sg13g2_fill_2 FILLER_28_40 ();
 sg13g2_fill_1 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_47 ();
 sg13g2_decap_8 FILLER_28_54 ();
 sg13g2_decap_8 FILLER_28_61 ();
 sg13g2_decap_8 FILLER_28_72 ();
 sg13g2_decap_8 FILLER_28_79 ();
 sg13g2_decap_8 FILLER_28_86 ();
 sg13g2_fill_2 FILLER_28_93 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_decap_4 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_106 ();
 sg13g2_decap_8 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_decap_4 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_fill_2 FILLER_28_153 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_25 ();
 sg13g2_fill_2 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_62 ();
 sg13g2_decap_8 FILLER_29_68 ();
 sg13g2_decap_4 FILLER_29_75 ();
 sg13g2_decap_8 FILLER_29_83 ();
 sg13g2_decap_4 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_fill_2 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_27 ();
 sg13g2_decap_8 FILLER_30_34 ();
 sg13g2_decap_8 FILLER_30_41 ();
 sg13g2_fill_2 FILLER_30_48 ();
 sg13g2_decap_8 FILLER_30_60 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_92 ();
 sg13g2_decap_8 FILLER_30_99 ();
 sg13g2_fill_2 FILLER_30_106 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_decap_4 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_139 ();
 sg13g2_decap_8 FILLER_30_146 ();
 sg13g2_decap_8 FILLER_30_153 ();
 sg13g2_decap_8 FILLER_30_160 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_decap_8 FILLER_31_120 ();
 sg13g2_decap_8 FILLER_31_127 ();
 sg13g2_decap_8 FILLER_31_134 ();
 sg13g2_decap_8 FILLER_31_141 ();
 sg13g2_fill_2 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_decap_4 FILLER_31_161 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_176 ();
 sg13g2_decap_4 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_47 ();
 sg13g2_decap_8 FILLER_32_54 ();
 sg13g2_decap_8 FILLER_32_61 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_decap_8 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_80 ();
 sg13g2_decap_4 FILLER_32_87 ();
 sg13g2_fill_1 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_decap_8 FILLER_32_149 ();
 sg13g2_decap_8 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_decap_8 FILLER_33_85 ();
 sg13g2_decap_8 FILLER_33_92 ();
 sg13g2_decap_8 FILLER_33_99 ();
 sg13g2_decap_4 FILLER_33_106 ();
 sg13g2_fill_2 FILLER_33_110 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_fill_1 FILLER_33_120 ();
 sg13g2_decap_8 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_decap_8 FILLER_33_155 ();
 sg13g2_decap_8 FILLER_33_162 ();
 sg13g2_decap_8 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_176 ();
 sg13g2_decap_4 FILLER_33_183 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_11 ();
 sg13g2_decap_8 FILLER_34_27 ();
 sg13g2_fill_1 FILLER_34_34 ();
 sg13g2_decap_4 FILLER_34_50 ();
 sg13g2_decap_4 FILLER_34_87 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_116 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_158 ();
 sg13g2_decap_8 FILLER_34_165 ();
 sg13g2_decap_8 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_179 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_4 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_2 FILLER_35_55 ();
 sg13g2_decap_8 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_79 ();
 sg13g2_decap_8 FILLER_35_86 ();
 sg13g2_decap_8 FILLER_35_93 ();
 sg13g2_decap_8 FILLER_35_100 ();
 sg13g2_decap_8 FILLER_35_107 ();
 sg13g2_fill_2 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_116 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_143 ();
 sg13g2_decap_8 FILLER_35_164 ();
 sg13g2_fill_1 FILLER_35_171 ();
 sg13g2_decap_4 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_186 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_31 ();
 sg13g2_fill_1 FILLER_36_39 ();
 sg13g2_fill_2 FILLER_36_43 ();
 sg13g2_decap_8 FILLER_36_48 ();
 sg13g2_decap_8 FILLER_36_65 ();
 sg13g2_decap_8 FILLER_36_72 ();
 sg13g2_decap_4 FILLER_36_79 ();
 sg13g2_fill_1 FILLER_36_83 ();
 sg13g2_fill_2 FILLER_36_103 ();
 sg13g2_decap_4 FILLER_36_118 ();
 sg13g2_fill_2 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_150 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_decap_4 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_fill_2 FILLER_37_55 ();
 sg13g2_fill_1 FILLER_37_57 ();
 sg13g2_decap_4 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_115 ();
 sg13g2_decap_8 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_fill_2 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_38 ();
 sg13g2_decap_8 FILLER_38_43 ();
 sg13g2_decap_8 FILLER_38_50 ();
 sg13g2_decap_8 FILLER_38_57 ();
 sg13g2_decap_8 FILLER_38_64 ();
 sg13g2_decap_8 FILLER_38_71 ();
 sg13g2_decap_4 FILLER_38_78 ();
 sg13g2_fill_1 FILLER_38_82 ();
 sg13g2_decap_4 FILLER_38_86 ();
 sg13g2_decap_4 FILLER_38_94 ();
 sg13g2_fill_2 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_106 ();
 sg13g2_decap_4 FILLER_38_113 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_decap_8 FILLER_38_125 ();
 sg13g2_decap_8 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_139 ();
 sg13g2_decap_8 FILLER_38_146 ();
 sg13g2_decap_8 FILLER_38_153 ();
 sg13g2_decap_8 FILLER_38_160 ();
 sg13g2_decap_8 FILLER_38_167 ();
 sg13g2_decap_8 FILLER_38_174 ();
 sg13g2_decap_8 FILLER_38_181 ();
 assign spine_bot_iw[1] = \genblk2[0].ctrl_ena_buf_I.z ;
 assign spine_bot_iw[11] = \genblk2[0].pad_ui_in_buf_I[0].z ;
 assign spine_bot_iw[12] = \genblk2[0].pad_ui_in_buf_I[1].z ;
 assign spine_bot_iw[13] = \genblk2[0].pad_ui_in_buf_I[2].z ;
 assign spine_bot_iw[14] = \genblk2[0].pad_ui_in_buf_I[3].z ;
 assign spine_bot_iw[15] = \genblk2[0].pad_ui_in_buf_I[4].z ;
 assign spine_bot_iw[16] = \genblk2[0].pad_ui_in_buf_I[5].z ;
 assign spine_bot_iw[17] = \genblk2[0].pad_ui_in_buf_I[6].z ;
 assign spine_bot_iw[18] = \genblk2[0].pad_ui_in_buf_I[7].z ;
 assign spine_bot_iw[19] = \genblk2[0].pad_ui_in_buf_I[8].z ;
 assign spine_bot_iw[20] = \genblk2[0].pad_ui_in_buf_I[9].z ;
 assign spine_bot_iw[21] = \genblk2[0].pad_uio_in_buf_I[0].z ;
 assign spine_bot_iw[22] = \genblk2[0].pad_uio_in_buf_I[1].z ;
 assign spine_bot_iw[23] = \genblk2[0].pad_uio_in_buf_I[2].z ;
 assign spine_bot_iw[24] = \genblk2[0].pad_uio_in_buf_I[3].z ;
 assign spine_bot_iw[25] = \genblk2[0].pad_uio_in_buf_I[4].z ;
 assign spine_bot_iw[26] = \genblk2[0].pad_uio_in_buf_I[5].z ;
 assign spine_bot_iw[27] = \genblk2[0].pad_uio_in_buf_I[6].z ;
 assign spine_bot_iw[28] = \genblk2[0].pad_uio_in_buf_I[7].z ;
 assign spine_bot_iw[2] = \genblk2[0].sel_cnt_buf_I[0].z ;
 assign spine_bot_iw[3] = \genblk2[0].sel_cnt_buf_I[1].z ;
 assign spine_bot_iw[4] = \genblk2[0].sel_cnt_buf_I[2].z ;
 assign spine_bot_iw[5] = \genblk2[0].sel_cnt_buf_I[3].z ;
 assign spine_bot_iw[6] = \genblk2[0].sel_cnt_buf_I[4].z ;
 assign spine_bot_iw[7] = \genblk2[0].sel_cnt_buf_I[5].z ;
 assign spine_bot_iw[8] = \genblk2[0].sel_cnt_buf_I[6].z ;
 assign spine_bot_iw[9] = \genblk2[0].sel_cnt_buf_I[7].z ;
 assign spine_bot_iw[10] = \genblk2[0].sel_cnt_buf_I[8].z ;
 assign spine_bot_iw[0] = \genblk2[0].tie_guard_I[0].lo ;
 assign spine_bot_iw[29] = \genblk2[0].tie_guard_I[1].lo ;
 assign spine_top_iw[1] = \genblk2[1].ctrl_ena_buf_I.z ;
 assign spine_top_iw[11] = \genblk2[1].pad_ui_in_buf_I[0].z ;
 assign spine_top_iw[12] = \genblk2[1].pad_ui_in_buf_I[1].z ;
 assign spine_top_iw[13] = \genblk2[1].pad_ui_in_buf_I[2].z ;
 assign spine_top_iw[14] = \genblk2[1].pad_ui_in_buf_I[3].z ;
 assign spine_top_iw[15] = \genblk2[1].pad_ui_in_buf_I[4].z ;
 assign spine_top_iw[16] = \genblk2[1].pad_ui_in_buf_I[5].z ;
 assign spine_top_iw[17] = \genblk2[1].pad_ui_in_buf_I[6].z ;
 assign spine_top_iw[18] = \genblk2[1].pad_ui_in_buf_I[7].z ;
 assign spine_top_iw[19] = \genblk2[1].pad_ui_in_buf_I[8].z ;
 assign spine_top_iw[20] = \genblk2[1].pad_ui_in_buf_I[9].z ;
 assign spine_top_iw[21] = \genblk2[1].pad_uio_in_buf_I[0].z ;
 assign spine_top_iw[22] = \genblk2[1].pad_uio_in_buf_I[1].z ;
 assign spine_top_iw[23] = \genblk2[1].pad_uio_in_buf_I[2].z ;
 assign spine_top_iw[24] = \genblk2[1].pad_uio_in_buf_I[3].z ;
 assign spine_top_iw[25] = \genblk2[1].pad_uio_in_buf_I[4].z ;
 assign spine_top_iw[26] = \genblk2[1].pad_uio_in_buf_I[5].z ;
 assign spine_top_iw[27] = \genblk2[1].pad_uio_in_buf_I[6].z ;
 assign spine_top_iw[28] = \genblk2[1].pad_uio_in_buf_I[7].z ;
 assign spine_top_iw[2] = \genblk2[1].sel_cnt_buf_I[0].z ;
 assign spine_top_iw[3] = \genblk2[1].sel_cnt_buf_I[1].z ;
 assign spine_top_iw[4] = \genblk2[1].sel_cnt_buf_I[2].z ;
 assign spine_top_iw[5] = \genblk2[1].sel_cnt_buf_I[3].z ;
 assign spine_top_iw[6] = \genblk2[1].sel_cnt_buf_I[4].z ;
 assign spine_top_iw[7] = \genblk2[1].sel_cnt_buf_I[5].z ;
 assign spine_top_iw[8] = \genblk2[1].sel_cnt_buf_I[6].z ;
 assign spine_top_iw[9] = \genblk2[1].sel_cnt_buf_I[7].z ;
 assign spine_top_iw[10] = \genblk2[1].sel_cnt_buf_I[8].z ;
 assign spine_top_iw[0] = \genblk2[1].tie_guard_I[0].lo ;
 assign spine_top_iw[29] = \genblk2[1].tie_guard_I[1].lo ;
 assign pad_uio_oex[0] = \uio_oe_obuf_I[0].z ;
 assign pad_uio_oex[1] = \uio_oe_obuf_I[1].z ;
 assign pad_uio_oex[2] = \uio_oe_obuf_I[2].z ;
 assign pad_uio_oex[3] = \uio_oe_obuf_I[3].z ;
 assign pad_uio_oex[4] = \uio_oe_obuf_I[4].z ;
 assign pad_uio_oex[5] = \uio_oe_obuf_I[5].z ;
 assign pad_uio_oex[6] = \uio_oe_obuf_I[6].z ;
 assign pad_uio_oex[7] = \uio_oe_obuf_I[7].z ;
 assign pad_uio_out[0] = \uio_out_obuf_I[0].z ;
 assign pad_uio_out[1] = \uio_out_obuf_I[1].z ;
 assign pad_uio_out[2] = \uio_out_obuf_I[2].z ;
 assign pad_uio_out[3] = \uio_out_obuf_I[3].z ;
 assign pad_uio_out[4] = \uio_out_obuf_I[4].z ;
 assign pad_uio_out[5] = \uio_out_obuf_I[5].z ;
 assign pad_uio_out[6] = \uio_out_obuf_I[6].z ;
 assign pad_uio_out[7] = \uio_out_obuf_I[7].z ;
 assign pad_uo_out[0] = \uo_out_obuf_I[0].z ;
 assign pad_uo_out[1] = \uo_out_obuf_I[1].z ;
 assign pad_uo_out[2] = \uo_out_obuf_I[2].z ;
 assign pad_uo_out[3] = \uo_out_obuf_I[3].z ;
 assign pad_uo_out[4] = \uo_out_obuf_I[4].z ;
 assign pad_uo_out[5] = \uo_out_obuf_I[5].z ;
 assign pad_uo_out[6] = \uo_out_obuf_I[6].z ;
 assign pad_uo_out[7] = \uo_out_obuf_I[7].z ;
endmodule
