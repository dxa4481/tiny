module tt_um_chip_rom (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire \addr_counter[0] ;
 wire \addr_counter[1] ;
 wire \addr_counter[2] ;
 wire \addr_counter[3] ;
 wire \addr_counter[4] ;
 wire \addr_counter[5] ;
 wire \addr_counter[6] ;
 wire \addr_counter[7] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire clknet_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net17;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net62;
 wire net63;
 wire net64;
 wire net65;

 sg13g2_inv_4 _183_ (.A(net61),
    .Y(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _184_ (.VDD(VPWR),
    .Y(_127_),
    .A(\addr_counter[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _185_ (.VDD(VPWR),
    .Y(_000_),
    .A(net33),
    .VSS(VGND));
 sg13g2_and2_1 _186_ (.A(net59),
    .B(net7),
    .X(_128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _187_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_128_),
    .Y(_129_),
    .A2(\addr_counter[6] ),
    .A1(_008_));
 sg13g2_a21o_2 _188_ (.A2(\addr_counter[6] ),
    .A1(_008_),
    .B1(_128_),
    .X(_130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _189_ (.A0(\addr_counter[5] ),
    .A1(net6),
    .S(net58),
    .X(_131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _190_ (.A(_129_),
    .B(net57),
    .Y(_132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _191_ (.Y(_133_),
    .A(net59),
    .B(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _192_ (.Y(_134_),
    .B(\addr_counter[0] ),
    .A_N(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _193_ (.A(_133_),
    .B(_134_),
    .X(_135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _194_ (.A0(\addr_counter[0] ),
    .A1(net1),
    .S(net59),
    .X(_136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _195_ (.A(net59),
    .B(\addr_counter[1] ),
    .Y(_137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _196_ (.A(net2),
    .B_N(net59),
    .Y(_138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _197_ (.A0(\addr_counter[1] ),
    .A1(net2),
    .S(net59),
    .X(_139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _198_ (.A(net55),
    .B(net52),
    .X(_140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _199_ (.Y(_141_),
    .A(net55),
    .B(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _200_ (.Y(_142_),
    .A(net3),
    .B(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _201_ (.Y(_143_),
    .B(\addr_counter[2] ),
    .A_N(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _202_ (.A0(\addr_counter[2] ),
    .A1(net3),
    .S(net59),
    .X(_144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _203_ (.Y(_145_),
    .B1(_142_),
    .B2(_143_),
    .A2(net52),
    .A1(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _204_ (.A(net48),
    .B_N(net54),
    .Y(_146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _205_ (.A(net49),
    .B_N(net52),
    .Y(_147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _206_ (.Y(_148_),
    .B(net50),
    .A_N(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _207_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net55),
    .A2(_147_),
    .Y(_149_),
    .B1(_145_));
 sg13g2_and2_1 _208_ (.A(net60),
    .B(net4),
    .X(_150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _209_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_150_),
    .Y(_151_),
    .A2(\addr_counter[3] ),
    .A1(_008_));
 sg13g2_mux2_1 _210_ (.A0(\addr_counter[3] ),
    .A1(net4),
    .S(net60),
    .X(_152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _211_ (.A(net58),
    .B(net5),
    .X(_153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _212_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_153_),
    .Y(_154_),
    .A2(\addr_counter[4] ),
    .A1(_008_));
 sg13g2_mux2_1 _213_ (.A0(\addr_counter[4] ),
    .A1(net5),
    .S(net58),
    .X(_155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _214_ (.A(_149_),
    .B(net46),
    .C(_154_),
    .Y(_156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _215_ (.A(net50),
    .B(net44),
    .X(_157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _216_ (.VDD(VPWR),
    .Y(_158_),
    .A(_157_),
    .VSS(VGND));
 sg13g2_nor2_1 _217_ (.A(net42),
    .B(_157_),
    .Y(_159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _218_ (.A(net55),
    .B(net52),
    .Y(_160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _219_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_161_),
    .B(net50),
    .A(net54));
 sg13g2_and2_1 _220_ (.A(net50),
    .B(net48),
    .X(_162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _221_ (.Y(_163_),
    .A(net52),
    .B(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _222_ (.A(net54),
    .B(_162_),
    .Y(_164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _223_ (.VDD(VPWR),
    .Y(_165_),
    .A(_164_),
    .VSS(VGND));
 sg13g2_xor2_1 _224_ (.B(_164_),
    .A(_159_),
    .X(_166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _225_ (.B1(_132_),
    .VDD(VPWR),
    .Y(_167_),
    .VSS(VGND),
    .A1(_156_),
    .A2(_166_));
 sg13g2_and2_1 _226_ (.A(_131_),
    .B(net43),
    .X(_168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _227_ (.Y(_169_),
    .A(net57),
    .B(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _228_ (.A(net55),
    .B(_137_),
    .C(_138_),
    .Y(_170_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net49));
 sg13g2_nand2_1 _229_ (.Y(_171_),
    .A(_151_),
    .B(_170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _230_ (.A(_145_),
    .B(_146_),
    .C(net46),
    .Y(_172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _231_ (.A(net54),
    .B(net48),
    .X(_173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _232_ (.A(_160_),
    .B(_173_),
    .Y(_174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _233_ (.B1(_171_),
    .VDD(VPWR),
    .Y(_175_),
    .VSS(VGND),
    .A1(_172_),
    .A2(_174_));
 sg13g2_nor2b_1 _234_ (.A(net50),
    .B_N(net48),
    .Y(_176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _235_ (.Y(_177_),
    .B(net49),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net52));
 sg13g2_nor2_2 _236_ (.A(net50),
    .B(net48),
    .Y(_178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _237_ (.A(net54),
    .B(net50),
    .C(net48),
    .Y(_179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _238_ (.A(_133_),
    .B(_134_),
    .C(net53),
    .D(net49),
    .X(_180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _239_ (.Y(_181_),
    .A(_135_),
    .B(_162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _240_ (.B1(_151_),
    .VDD(VPWR),
    .Y(_182_),
    .VSS(VGND),
    .A1(_179_),
    .A2(_180_));
 sg13g2_or4_1 _241_ (.A(_145_),
    .B(_146_),
    .C(_179_),
    .D(_180_),
    .X(_016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _242_ (.A(net42),
    .B_N(net57),
    .Y(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _243_ (.Y(_018_),
    .A(net57),
    .B(_154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _244_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_182_),
    .A2(_016_),
    .Y(_019_),
    .B1(_018_));
 sg13g2_or2_1 _245_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_020_),
    .B(net44),
    .A(net48));
 sg13g2_nor2_2 _246_ (.A(_131_),
    .B(net43),
    .Y(_021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _247_ (.B1(net46),
    .VDD(VPWR),
    .Y(_022_),
    .VSS(VGND),
    .A1(_140_),
    .A2(_179_));
 sg13g2_and2_1 _248_ (.A(_021_),
    .B(_022_),
    .X(_023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _249_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_023_),
    .C1(_019_),
    .B1(_020_),
    .A1(_168_),
    .Y(_024_),
    .A2(_175_));
 sg13g2_o21ai_1 _250_ (.B1(_167_),
    .VDD(VPWR),
    .Y(_025_),
    .VSS(VGND),
    .A1(_130_),
    .A2(_024_));
 sg13g2_and2_1 _251_ (.A(net60),
    .B(net8),
    .X(_026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _252_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_026_),
    .Y(_027_),
    .A2(\addr_counter[7] ),
    .A1(_008_));
 sg13g2_o21ai_1 _253_ (.B1(net45),
    .VDD(VPWR),
    .Y(_028_),
    .VSS(VGND),
    .A1(net51),
    .A2(net49));
 sg13g2_or3_1 _254_ (.A(_169_),
    .B(net41),
    .C(_028_),
    .X(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _255_ (.A(_129_),
    .B(_169_),
    .C(net41),
    .Y(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _256_ (.A(_129_),
    .B(_164_),
    .C(_029_),
    .Y(_031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _257_ (.A2(net41),
    .A1(_025_),
    .B1(_031_),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _258_ (.A(net44),
    .B_N(net54),
    .Y(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _259_ (.Y(_033_),
    .A(_178_),
    .B(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _260_ (.A(_018_),
    .B(_033_),
    .Y(_034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _261_ (.A(_129_),
    .B(_034_),
    .Y(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _262_ (.B1(_130_),
    .VDD(VPWR),
    .Y(_036_),
    .VSS(VGND),
    .A1(_018_),
    .A2(_033_));
 sg13g2_a21oi_1 _263_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net44),
    .A2(_162_),
    .Y(_037_),
    .B1(net42));
 sg13g2_o21ai_1 _264_ (.B1(_154_),
    .VDD(VPWR),
    .Y(_038_),
    .VSS(VGND),
    .A1(_151_),
    .A2(_163_));
 sg13g2_nor2_1 _265_ (.A(_160_),
    .B(_020_),
    .Y(_039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _266_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_157_),
    .A2(_173_),
    .Y(_040_),
    .B1(_039_));
 sg13g2_a221oi_1 _267_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net42),
    .C1(net57),
    .B1(_040_),
    .A1(_182_),
    .Y(_041_),
    .A2(_037_));
 sg13g2_nand2_1 _268_ (.Y(_042_),
    .A(_145_),
    .B(_161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _269_ (.B(net44),
    .C(_161_),
    .A(_145_),
    .Y(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _270_ (.B(_142_),
    .C(_143_),
    .A(_135_),
    .Y(_044_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net46));
 sg13g2_nand3_1 _271_ (.B(_177_),
    .C(_044_),
    .A(_141_),
    .Y(_045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _272_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net54),
    .A2(net48),
    .Y(_046_),
    .B1(net44));
 sg13g2_xnor2_1 _273_ (.Y(_047_),
    .A(net45),
    .B(_173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _274_ (.A(net51),
    .B(_169_),
    .Y(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _275_ (.A(_161_),
    .B(_020_),
    .Y(_049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _276_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_017_),
    .C1(_130_),
    .B1(_049_),
    .A1(_047_),
    .Y(_050_),
    .A2(_048_));
 sg13g2_o21ai_1 _277_ (.B1(_050_),
    .VDD(VPWR),
    .Y(_051_),
    .VSS(VGND),
    .A1(_018_),
    .A2(_043_));
 sg13g2_a21oi_1 _278_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_021_),
    .A2(_045_),
    .Y(_052_),
    .B1(_051_));
 sg13g2_o21ai_1 _279_ (.B1(net41),
    .VDD(VPWR),
    .Y(_053_),
    .VSS(VGND),
    .A1(_036_),
    .A2(_041_));
 sg13g2_nand2_1 _280_ (.Y(_054_),
    .A(net45),
    .B(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _281_ (.A(_054_),
    .B_N(net51),
    .Y(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _282_ (.B(net47),
    .C(_030_),
    .A(_147_),
    .Y(_056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _283_ (.B1(_056_),
    .VDD(VPWR),
    .Y(net10),
    .VSS(VGND),
    .A1(_052_),
    .A2(_053_));
 sg13g2_nor3_1 _284_ (.A(_162_),
    .B(_173_),
    .C(_178_),
    .Y(_057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _285_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_058_),
    .B(_057_),
    .A(_054_));
 sg13g2_o21ai_1 _286_ (.B1(_017_),
    .VDD(VPWR),
    .Y(_059_),
    .VSS(VGND),
    .A1(_180_),
    .A2(_028_));
 sg13g2_a21oi_1 _287_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net46),
    .A2(_160_),
    .Y(_060_),
    .B1(_140_));
 sg13g2_nand2_1 _288_ (.Y(_061_),
    .A(_168_),
    .B(_060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _289_ (.Y(_062_),
    .B1(_059_),
    .B2(_061_),
    .A2(_178_),
    .A1(_151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _290_ (.B1(net52),
    .VDD(VPWR),
    .Y(_063_),
    .VSS(VGND),
    .A1(net55),
    .A2(_144_));
 sg13g2_o21ai_1 _291_ (.B1(_063_),
    .VDD(VPWR),
    .Y(_064_),
    .VSS(VGND),
    .A1(_146_),
    .A2(_151_));
 sg13g2_a21o_1 _292_ (.A2(_064_),
    .A1(_021_),
    .B1(_130_),
    .X(_065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _293_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net46),
    .Y(_066_),
    .A2(net53),
    .A1(net56));
 sg13g2_nand2b_1 _294_ (.Y(_067_),
    .B(net43),
    .A_N(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _295_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_177_),
    .A2(_066_),
    .Y(_068_),
    .B1(_067_));
 sg13g2_o21ai_1 _296_ (.B1(_068_),
    .VDD(VPWR),
    .Y(_069_),
    .VSS(VGND),
    .A1(_149_),
    .A2(_151_));
 sg13g2_nor3_1 _297_ (.A(_157_),
    .B(_176_),
    .C(_032_),
    .Y(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _298_ (.B1(_021_),
    .VDD(VPWR),
    .Y(_071_),
    .VSS(VGND),
    .A1(_173_),
    .A2(_070_));
 sg13g2_a21oi_1 _299_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_017_),
    .A2(_049_),
    .Y(_072_),
    .B1(_129_));
 sg13g2_and3_1 _300_ (.X(_073_),
    .A(_069_),
    .B(_071_),
    .C(_072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _301_ (.B1(net41),
    .VDD(VPWR),
    .Y(_074_),
    .VSS(VGND),
    .A1(_062_),
    .A2(_065_));
 sg13g2_o21ai_1 _302_ (.B1(_058_),
    .VDD(VPWR),
    .Y(net11),
    .VSS(VGND),
    .A1(_073_),
    .A2(_074_));
 sg13g2_nor2_1 _303_ (.A(net44),
    .B(_178_),
    .Y(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _304_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_075_),
    .C1(_038_),
    .B1(_181_),
    .A1(net46),
    .Y(_076_),
    .A2(_160_));
 sg13g2_a221oi_1 _305_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_135_),
    .C1(_151_),
    .B1(_178_),
    .A1(_145_),
    .Y(_077_),
    .A2(_161_));
 sg13g2_nor3_1 _306_ (.A(_154_),
    .B(_172_),
    .C(_077_),
    .Y(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _307_ (.B1(_132_),
    .VDD(VPWR),
    .Y(_079_),
    .VSS(VGND),
    .A1(_076_),
    .A2(_078_));
 sg13g2_nand2_1 _308_ (.Y(_080_),
    .A(_042_),
    .B(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _309_ (.B1(_135_),
    .VDD(VPWR),
    .Y(_081_),
    .VSS(VGND),
    .A1(net51),
    .A2(net45));
 sg13g2_a21oi_1 _310_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_146_),
    .A2(_158_),
    .Y(_082_),
    .B1(_169_));
 sg13g2_a21oi_1 _311_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_147_),
    .A2(net46),
    .Y(_083_),
    .B1(_130_));
 sg13g2_nand2_1 _312_ (.Y(_084_),
    .A(_148_),
    .B(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _313_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_083_),
    .A2(_084_),
    .Y(_085_),
    .B1(_018_));
 sg13g2_a221oi_1 _314_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_082_),
    .C1(_085_),
    .B1(_081_),
    .A1(_023_),
    .Y(_086_),
    .A2(_080_));
 sg13g2_o21ai_1 _315_ (.B1(_079_),
    .VDD(VPWR),
    .Y(_087_),
    .VSS(VGND),
    .A1(_035_),
    .A2(_086_));
 sg13g2_a21o_1 _316_ (.A2(_087_),
    .A1(net41),
    .B1(_055_),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _317_ (.B(_177_),
    .C(_030_),
    .A(net47),
    .Y(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _318_ (.A(_131_),
    .B(_170_),
    .C(_066_),
    .Y(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _319_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_020_),
    .A2(_089_),
    .Y(_090_),
    .B1(_021_));
 sg13g2_a22oi_1 _320_ (.Y(_091_),
    .B1(_177_),
    .B2(_066_),
    .A2(_163_),
    .A1(_161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _321_ (.A(_140_),
    .B(_160_),
    .C(_020_),
    .Y(_092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _322_ (.A(net43),
    .B(_091_),
    .C(_092_),
    .Y(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _323_ (.B1(_072_),
    .VDD(VPWR),
    .Y(_094_),
    .VSS(VGND),
    .A1(_090_),
    .A2(_093_));
 sg13g2_nand2_1 _324_ (.Y(_095_),
    .A(_141_),
    .B(_148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _325_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net45),
    .C1(_018_),
    .B1(_095_),
    .A1(_165_),
    .Y(_096_),
    .A2(_066_));
 sg13g2_a221oi_1 _326_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_135_),
    .C1(_169_),
    .B1(_028_),
    .A1(net45),
    .Y(_097_),
    .A2(_173_));
 sg13g2_nor4_1 _327_ (.A(_130_),
    .B(_023_),
    .C(_096_),
    .D(_097_),
    .Y(_098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _328_ (.Y(_099_),
    .A(_027_),
    .B(_094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _329_ (.B1(_088_),
    .VDD(VPWR),
    .Y(net13),
    .VSS(VGND),
    .A1(_098_),
    .A2(_099_));
 sg13g2_o21ai_1 _330_ (.B1(net57),
    .VDD(VPWR),
    .Y(_100_),
    .VSS(VGND),
    .A1(_161_),
    .A2(_020_));
 sg13g2_a22oi_1 _331_ (.Y(_101_),
    .B1(_176_),
    .B2(_032_),
    .A2(_157_),
    .A1(_146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _332_ (.Y(_102_),
    .A(_154_),
    .B(_101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _333_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_100_),
    .A2(_102_),
    .Y(_103_),
    .B1(_130_));
 sg13g2_nand3_1 _334_ (.B(_178_),
    .C(_032_),
    .A(net42),
    .Y(_104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _335_ (.B(_169_),
    .C(_100_),
    .A(_130_),
    .Y(_105_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_104_));
 sg13g2_nand2b_1 _336_ (.Y(_106_),
    .B(_105_),
    .A_N(_103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _337_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net56),
    .A2(_162_),
    .Y(_107_),
    .B1(_029_));
 sg13g2_mux2_1 _338_ (.A0(_107_),
    .A1(net41),
    .S(_106_),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _339_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net55),
    .A2(_147_),
    .Y(_108_),
    .B1(_088_));
 sg13g2_nor3_1 _340_ (.A(_162_),
    .B(_179_),
    .C(_046_),
    .Y(_109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _341_ (.B1(net42),
    .VDD(VPWR),
    .Y(_110_),
    .VSS(VGND),
    .A1(_049_),
    .A2(_109_));
 sg13g2_nand2_1 _342_ (.Y(_111_),
    .A(_162_),
    .B(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _343_ (.A2(_111_),
    .A1(_043_),
    .B1(net42),
    .X(_112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _344_ (.B(net57),
    .C(_110_),
    .A(_129_),
    .Y(_113_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_112_));
 sg13g2_nand3b_1 _345_ (.B(net44),
    .C(net54),
    .Y(_114_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net50));
 sg13g2_or2_1 _346_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_115_),
    .B(_170_),
    .A(_151_));
 sg13g2_a21oi_1 _347_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_178_),
    .A2(_032_),
    .Y(_116_),
    .B1(_154_));
 sg13g2_a22oi_1 _348_ (.Y(_117_),
    .B1(_115_),
    .B2(_116_),
    .A2(_114_),
    .A1(_037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _349_ (.Y(_118_),
    .B(_132_),
    .A_N(_117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _350_ (.B(_021_),
    .C(_083_),
    .Y(_119_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_170_));
 sg13g2_nand3_1 _351_ (.B(_118_),
    .C(_119_),
    .A(_113_),
    .Y(_120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _352_ (.A2(_120_),
    .A1(net41),
    .B1(_108_),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _353_ (.A(_054_),
    .B_N(_095_),
    .Y(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _354_ (.B(net34),
    .A(net33),
    .X(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _355_ (.B(net33),
    .C(net34),
    .A(net64),
    .Y(_121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _356_ (.A2(net34),
    .A1(net33),
    .B1(net64),
    .X(_122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _357_ (.A(_121_),
    .B(_122_),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _358_ (.A(_127_),
    .B(_121_),
    .Y(_123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _359_ (.Y(_003_),
    .A(net62),
    .B(_121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _360_ (.A(net39),
    .B(_123_),
    .X(_124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _361_ (.B(_123_),
    .A(net39),
    .X(_004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _362_ (.B(_124_),
    .A(net37),
    .X(_005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _363_ (.B(net65),
    .C(_124_),
    .A(net37),
    .Y(_125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _364_ (.A2(_124_),
    .A1(net37),
    .B1(net65),
    .X(_126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _365_ (.A(_125_),
    .B(_126_),
    .X(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _366_ (.Y(_007_),
    .A(net35),
    .B(_125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _367_ (.VDD(VPWR),
    .Y(_009_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _368_ (.VDD(VPWR),
    .Y(_010_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _369_ (.VDD(VPWR),
    .Y(_011_),
    .A(net58),
    .VSS(VGND));
 sg13g2_inv_1 _370_ (.VDD(VPWR),
    .Y(_012_),
    .A(net58),
    .VSS(VGND));
 sg13g2_inv_1 _371_ (.VDD(VPWR),
    .Y(_013_),
    .A(net58),
    .VSS(VGND));
 sg13g2_inv_1 _372_ (.VDD(VPWR),
    .Y(_014_),
    .A(net58),
    .VSS(VGND));
 sg13g2_inv_1 _373_ (.VDD(VPWR),
    .Y(_015_),
    .A(net58),
    .VSS(VGND));
 sg13g2_dfrbpq_2 _374_ (.RESET_B(_008_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_000_),
    .Q(\addr_counter[0] ),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _375_ (.RESET_B(_009_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_001_),
    .Q(\addr_counter[1] ),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _376_ (.RESET_B(_010_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_002_),
    .Q(\addr_counter[2] ),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _377_ (.RESET_B(_011_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net63),
    .Q(\addr_counter[3] ),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _378_ (.RESET_B(_012_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net40),
    .Q(\addr_counter[4] ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _379_ (.RESET_B(_013_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net38),
    .Q(\addr_counter[5] ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _380_ (.RESET_B(_014_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_006_),
    .Q(\addr_counter[6] ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _381_ (.RESET_B(_015_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net36),
    .Q(\addr_counter[7] ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_chip_rom_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net18));
 sg13g2_tielo tt_um_chip_rom_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net19));
 sg13g2_tielo tt_um_chip_rom_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net20));
 sg13g2_tielo tt_um_chip_rom_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net21));
 sg13g2_tielo tt_um_chip_rom_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net22));
 sg13g2_tielo tt_um_chip_rom_23 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net23));
 sg13g2_tielo tt_um_chip_rom_24 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net24));
 sg13g2_tielo tt_um_chip_rom_25 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net25));
 sg13g2_tielo tt_um_chip_rom_26 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net26));
 sg13g2_tielo tt_um_chip_rom_27 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net27));
 sg13g2_tielo tt_um_chip_rom_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net28));
 sg13g2_tielo tt_um_chip_rom_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net29));
 sg13g2_tielo tt_um_chip_rom_30 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net30));
 sg13g2_tielo tt_um_chip_rom_31 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net31));
 sg13g2_tielo tt_um_chip_rom_32 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net32));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout41 (.A(_027_),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout42 (.A(_155_),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout43 (.A(_155_),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout44 (.A(net47),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout45 (.A(net47),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout46 (.A(net47),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout47 (.A(_152_),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout48 (.A(net49),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout49 (.A(_144_),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout50 (.A(net53),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout51 (.A(net53),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout52 (.A(net53),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout53 (.A(_139_),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout54 (.A(net56),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout55 (.A(net56),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout56 (.A(_136_),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout57 (.A(_131_),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout58 (.A(net61),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout59 (.A(net60),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout60 (.A(net61),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout61 (.A(rst_n),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo tt_um_chip_rom_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net17));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\addr_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold2 (.A(\addr_counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold3 (.A(\addr_counter[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold4 (.A(_007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold5 (.A(\addr_counter[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold6 (.A(_005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold7 (.A(\addr_counter[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold8 (.A(_004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold9 (.A(\addr_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold10 (.A(_003_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold11 (.A(\addr_counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold12 (.A(\addr_counter[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net65));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_407 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule
