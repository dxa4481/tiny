module tt_ihp_wrapper (iovdd,
    iovss,
    vgnd,
    vdpwr,
    pad_raw);
 inout iovdd;
 inout iovss;
 inout vgnd;
 inout vdpwr;
 inout [63:0] pad_raw;

 wire \gpio[0].gpio_I.pad_ana ;
 wire \gpio[0].gpio_I.pad_in ;
 wire \gpio[0].gpio_I.pad_oe ;
 wire \gpio[10].gpio_I.pad_ana ;
 wire \gpio[10].gpio_I.pad_in ;
 wire \gpio[10].gpio_I.pad_out ;
 wire \gpio[11].gpio_I.pad_ana ;
 wire \gpio[11].gpio_I.pad_in ;
 wire \gpio[11].gpio_I.pad_out ;
 wire \gpio[12].gpio_I.pad_ana ;
 wire \gpio[12].gpio_I.pad_in ;
 wire \gpio[12].gpio_I.pad_out ;
 wire \gpio[13].gpio_I.pad_ana ;
 wire \gpio[13].gpio_I.pad_in ;
 wire \gpio[13].gpio_I.pad_out ;
 wire \gpio[14].gpio_I.pad_ana ;
 wire \gpio[14].gpio_I.pad_in ;
 wire \gpio[14].gpio_I.pad_out ;
 wire \gpio[15].gpio_I.pad_ana ;
 wire \gpio[15].gpio_I.pad_in ;
 wire \gpio[15].gpio_I.pad_out ;
 wire \gpio[18].gpio_I.pad_ana ;
 wire \gpio[18].gpio_I.pad_in ;
 wire \gpio[18].gpio_I.pad_oe ;
 wire \gpio[19].gpio_I.pad_ana ;
 wire \gpio[19].gpio_I.pad_in ;
 wire \gpio[1].gpio_I.pad_ana ;
 wire \gpio[1].gpio_I.pad_in ;
 wire \gpio[20].gpio_I.pad_ana ;
 wire \gpio[20].gpio_I.pad_in ;
 wire \gpio[21].gpio_I.pad_ana ;
 wire \gpio[21].gpio_I.pad_in ;
 wire \gpio[24].gpio_I.pad_ana ;
 wire \gpio[24].gpio_I.pad_in ;
 wire \gpio[25].gpio_I.pad_ana ;
 wire \gpio[25].gpio_I.pad_in ;
 wire \gpio[26].gpio_I.pad_ana ;
 wire \gpio[26].gpio_I.pad_in ;
 wire \gpio[27].gpio_I.pad_ana ;
 wire \gpio[27].gpio_I.pad_in ;
 wire \gpio[2].gpio_I.pad_ana ;
 wire \gpio[2].gpio_I.pad_in ;
 wire \gpio[32].gpio_I.pad_ana ;
 wire \gpio[32].gpio_I.pad_in ;
 wire \gpio[32].gpio_I.pad_oe ;
 wire \gpio[32].gpio_I.pad_out ;
 wire \gpio[33].gpio_I.pad_ana ;
 wire \gpio[33].gpio_I.pad_in ;
 wire \gpio[33].gpio_I.pad_oe ;
 wire \gpio[33].gpio_I.pad_out ;
 wire \gpio[34].gpio_I.pad_ana ;
 wire \gpio[34].gpio_I.pad_in ;
 wire \gpio[34].gpio_I.pad_oe ;
 wire \gpio[34].gpio_I.pad_out ;
 wire \gpio[35].gpio_I.pad_ana ;
 wire \gpio[35].gpio_I.pad_in ;
 wire \gpio[35].gpio_I.pad_oe ;
 wire \gpio[35].gpio_I.pad_out ;
 wire \gpio[36].gpio_I.pad_ana ;
 wire \gpio[36].gpio_I.pad_in ;
 wire \gpio[36].gpio_I.pad_oe ;
 wire \gpio[36].gpio_I.pad_out ;
 wire \gpio[37].gpio_I.pad_ana ;
 wire \gpio[37].gpio_I.pad_in ;
 wire \gpio[37].gpio_I.pad_oe ;
 wire \gpio[37].gpio_I.pad_out ;
 wire \gpio[38].gpio_I.pad_ana ;
 wire \gpio[38].gpio_I.pad_in ;
 wire \gpio[38].gpio_I.pad_oe ;
 wire \gpio[38].gpio_I.pad_out ;
 wire \gpio[39].gpio_I.pad_ana ;
 wire \gpio[39].gpio_I.pad_in ;
 wire \gpio[39].gpio_I.pad_oe ;
 wire \gpio[39].gpio_I.pad_out ;
 wire \gpio[3].gpio_I.pad_ana ;
 wire \gpio[3].gpio_I.pad_in ;
 wire \gpio[40].gpio_I.pad_ana ;
 wire \gpio[40].gpio_I.pad_in ;
 wire \gpio[41].gpio_I.pad_ana ;
 wire \gpio[41].gpio_I.pad_in ;
 wire \gpio[42].gpio_I.pad_ana ;
 wire \gpio[42].gpio_I.pad_in ;
 wire \gpio[43].gpio_I.pad_ana ;
 wire \gpio[43].gpio_I.pad_in ;
 wire \gpio[44].gpio_I.pad_ana ;
 wire \gpio[44].gpio_I.pad_in ;
 wire \gpio[45].gpio_I.pad_ana ;
 wire \gpio[45].gpio_I.pad_in ;
 wire \gpio[46].gpio_I.pad_ana ;
 wire \gpio[46].gpio_I.pad_in ;
 wire \gpio[47].gpio_I.pad_ana ;
 wire \gpio[47].gpio_I.pad_in ;
 wire \gpio[48].gpio_I.pad_ana ;
 wire \gpio[48].gpio_I.pad_in ;
 wire \gpio[49].gpio_I.pad_ana ;
 wire \gpio[49].gpio_I.pad_in ;
 wire \gpio[4].gpio_I.pad_ana ;
 wire \gpio[4].gpio_I.pad_in ;
 wire \gpio[52].gpio_I.pad_ana ;
 wire \gpio[52].gpio_I.pad_in ;
 wire \gpio[53].gpio_I.pad_ana ;
 wire \gpio[53].gpio_I.pad_in ;
 wire \gpio[54].gpio_I.pad_ana ;
 wire \gpio[54].gpio_I.pad_in ;
 wire \gpio[55].gpio_I.pad_ana ;
 wire \gpio[55].gpio_I.pad_in ;
 wire \gpio[58].gpio_I.pad_ana ;
 wire \gpio[58].gpio_I.pad_in ;
 wire \gpio[59].gpio_I.pad_ana ;
 wire \gpio[59].gpio_I.pad_in ;
 wire \gpio[5].gpio_I.pad_ana ;
 wire \gpio[5].gpio_I.pad_in ;
 wire \gpio[60].gpio_I.pad_ana ;
 wire \gpio[60].gpio_I.pad_in ;
 wire \gpio[61].gpio_I.pad_ana ;
 wire \gpio[61].gpio_I.pad_in ;
 wire \gpio[8].gpio_I.pad_ana ;
 wire \gpio[8].gpio_I.pad_in ;
 wire \gpio[8].gpio_I.pad_out ;
 wire \gpio[9].gpio_I.pad_ana ;
 wire \gpio[9].gpio_I.pad_in ;
 wire \gpio[9].gpio_I.pad_out ;
 wire \top_I.branch[0].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.l_addr[0] ;
 wire \top_I.branch[0].check_mask.l_k_one ;
 wire \top_I.branch[0].check_mask.l_spine_iw[0] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[10] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[11] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[12] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[13] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[14] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[15] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[16] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[17] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[18] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[19] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[1] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[20] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[21] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[22] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[23] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[24] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[25] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[26] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[27] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[28] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[29] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[2] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[3] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[4] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[5] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[6] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[7] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[8] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[9] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[0] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[10] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[11] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[12] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[13] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[14] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[15] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[16] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[17] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[18] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[19] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[1] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[20] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[21] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[22] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[23] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[24] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[25] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[2] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[3] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[4] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[5] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[6] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[7] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[8] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[9] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.l_addr[0] ;
 wire \top_I.branch[10].check_mask.l_addr[1] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.l_addr[0] ;
 wire \top_I.branch[13].check_mask.l_addr[1] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[0] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[10] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[11] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[12] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[13] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[14] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[15] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[16] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[17] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[18] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[19] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[1] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[20] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[21] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[22] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[23] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[24] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[25] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[26] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[27] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[28] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[29] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[2] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[3] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[4] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[5] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[6] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[7] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[8] ;
 wire \top_I.branch[13].check_mask.l_spine_iw[9] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[0] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[10] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[11] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[12] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[13] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[14] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[15] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[16] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[17] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[18] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[19] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[1] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[20] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[21] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[22] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[23] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[24] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[25] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[2] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[3] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[4] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[5] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[6] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[7] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[8] ;
 wire \top_I.branch[13].check_mask.l_spine_ow[9] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.l_addr[0] ;
 wire \top_I.branch[14].check_mask.l_addr[3] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.l_addr[0] ;
 wire \top_I.branch[15].check_mask.l_addr[3] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.l_addr[0] ;
 wire \top_I.branch[16].check_mask.l_addr[3] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.l_addr[0] ;
 wire \top_I.branch[17].check_mask.l_addr[3] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.l_addr[0] ;
 wire \top_I.branch[18].check_mask.l_addr[1] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.l_addr[0] ;
 wire \top_I.branch[19].check_mask.l_addr[1] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.l_addr[0] ;
 wire \top_I.branch[1].check_mask.l_k_one ;
 wire \top_I.branch[2].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.l_addr[0] ;
 wire \top_I.branch[2].check_mask.l_addr[1] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.l_addr[0] ;
 wire \top_I.branch[3].check_mask.l_addr[1] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.l_addr[0] ;
 wire \top_I.branch[4].check_mask.l_addr[1] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.l_addr[0] ;
 wire \top_I.branch[5].check_mask.l_addr[1] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.l_addr[0] ;
 wire \top_I.branch[7].check_mask.l_addr[2] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.l_addr[0] ;
 wire \top_I.branch[8].check_mask.l_addr[2] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.l_addr[0] ;
 wire \top_I.branch[9].check_mask.l_addr[2] ;
 wire vapwr;
 wire \top_I.branch[0].check_mask.block[0].um_I.block_0_0.vdpwr ;
 wire \top_I.branch[0].check_mask.block[1].um_I.block_0_1.vdpwr ;
 wire \top_I.branch[10].check_mask.block[0].um_I.block_10_0.vdpwr ;
 wire \top_I.branch[10].check_mask.block[2].um_I.block_10_2.vdpwr ;
 wire \top_I.branch[16].check_mask.block[11].um_I.block_16_11.vdpwr ;
 wire \top_I.branch[16].check_mask.block[1].um_I.block_16_1.vdpwr ;
 wire \top_I.branch[16].check_mask.block[3].um_I.block_16_3.vdpwr ;
 wire \top_I.branch[16].check_mask.block[5].um_I.block_16_5.vdpwr ;
 wire \top_I.branch[16].check_mask.block[7].um_I.block_16_7.vdpwr ;
 wire \top_I.branch[16].check_mask.block[9].um_I.block_16_9.vdpwr ;

 sg13g2_IOPadIn \gpio[0].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[0].gpio_I.pad_in ),
    .pad(pad_raw[0]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut30mA \gpio[10].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[10].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[10]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut30mA \gpio[11].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[11].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[11]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut30mA \gpio[12].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[12].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[12]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut30mA \gpio[13].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[13].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[13]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut30mA \gpio[14].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[14].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[14]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut30mA \gpio[15].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[15].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[15]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[16].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[17].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[18].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[19].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[1].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[1].gpio_I.pad_in ),
    .pad(pad_raw[1]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[20].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[21].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[22].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[23].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[24].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[25].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[26].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[27].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadVss \gpio[28].gpio_I.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadVdd \gpio[29].gpio_I.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[2].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[2].gpio_I.pad_in ),
    .pad(pad_raw[2]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[30].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[31].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut30mA \gpio[32].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[32].gpio_I.pad_out ),
    .c2p_en(\gpio[32].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[32].gpio_I.pad_in ),
    .pad(pad_raw[32]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut30mA \gpio[33].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[33].gpio_I.pad_out ),
    .c2p_en(\gpio[33].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[33].gpio_I.pad_in ),
    .pad(pad_raw[33]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut30mA \gpio[34].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[34].gpio_I.pad_out ),
    .c2p_en(\gpio[34].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[34].gpio_I.pad_in ),
    .pad(pad_raw[34]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut30mA \gpio[35].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[35].gpio_I.pad_out ),
    .c2p_en(\gpio[35].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[35].gpio_I.pad_in ),
    .pad(pad_raw[35]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut30mA \gpio[36].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[36].gpio_I.pad_out ),
    .c2p_en(\gpio[36].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[36].gpio_I.pad_in ),
    .pad(pad_raw[36]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut30mA \gpio[37].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[37].gpio_I.pad_out ),
    .c2p_en(\gpio[37].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[37].gpio_I.pad_in ),
    .pad(pad_raw[37]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut30mA \gpio[38].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[38].gpio_I.pad_out ),
    .c2p_en(\gpio[38].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[38].gpio_I.pad_in ),
    .pad(pad_raw[38]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut30mA \gpio[39].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[39].gpio_I.pad_out ),
    .c2p_en(\gpio[39].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[39].gpio_I.pad_in ),
    .pad(pad_raw[39]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[3].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[3].gpio_I.pad_in ),
    .pad(pad_raw[3]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[40].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[40].gpio_I.pad_in ),
    .pad(pad_raw[40]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[41].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[41].gpio_I.pad_in ),
    .pad(pad_raw[41]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[42].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[42].gpio_I.pad_in ),
    .pad(pad_raw[42]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[43].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[43].gpio_I.pad_in ),
    .pad(pad_raw[43]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[44].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[44].gpio_I.pad_in ),
    .pad(pad_raw[44]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[45].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[45].gpio_I.pad_in ),
    .pad(pad_raw[45]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[46].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[46].gpio_I.pad_in ),
    .pad(pad_raw[46]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[47].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[47].gpio_I.pad_in ),
    .pad(pad_raw[47]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[48].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[48].gpio_I.pad_in ),
    .pad(pad_raw[48]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[49].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[49].gpio_I.pad_in ),
    .pad(pad_raw[49]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[4].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[4].gpio_I.pad_in ),
    .pad(pad_raw[4]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[50].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[51].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[52].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[53].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[54].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[55].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[56].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[57].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[58].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[59].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[5].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[5].gpio_I.pad_in ),
    .pad(pad_raw[5]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[60].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[61].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadVss \gpio[62].gpio_I.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadVdd \gpio[63].gpio_I.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[6].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[7].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut30mA \gpio[8].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[8].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[8]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut30mA \gpio[9].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.c2p(\gpio[9].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[9]),
    .vdd(vdpwr),
    .vss(vgnd));
 tt_pg_1v5_ll_1 \top_I.branch[0].check_mask.block[0].um_I.block_0_0.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[0].check_mask.block[0].um_I.block_0_0.vdpwr ),
    .ctrl(\top_I.branch[0].check_mask.block[0].um_I.pg_ena ));
 tt_um_chip_rom \top_I.branch[0].check_mask.block[0].um_I.block_0_0.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[0].check_mask.block[0].um_I.block_0_0.vdpwr ),
    .clk(\top_I.branch[0].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[0] }));
 tt_pg_1v5_ll_1 \top_I.branch[0].check_mask.block[1].um_I.block_0_1.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[0].check_mask.block[1].um_I.block_0_1.vdpwr ),
    .ctrl(\top_I.branch[0].check_mask.block[1].um_I.pg_ena ));
 tt_um_factory_test \top_I.branch[0].check_mask.block[1].um_I.block_0_1.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[0].check_mask.block[1].um_I.block_0_1.vdpwr ),
    .clk(\top_I.branch[0].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[0] }));
 tt_mux \top_I.branch[0].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[0].check_mask.l_k_one ),
    .k_zero(\top_I.branch[0].check_mask.l_addr[0] ),
    .addr({\top_I.branch[0].check_mask.l_addr[0] ,
    \top_I.branch[0].check_mask.l_addr[0] ,
    \top_I.branch[0].check_mask.l_addr[0] ,
    \top_I.branch[0].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[0].check_mask.block[11].um_I.ena ,
    \top_I.branch[0].check_mask.block[10].um_I.ena ,
    \top_I.branch[0].check_mask.block[9].um_I.ena ,
    \top_I.branch[0].check_mask.block[8].um_I.ena ,
    \top_I.branch[0].check_mask.block[7].um_I.ena ,
    \top_I.branch[0].check_mask.block[6].um_I.ena ,
    \top_I.branch[0].check_mask.block[5].um_I.ena ,
    \top_I.branch[0].check_mask.block[4].um_I.ena ,
    \top_I.branch[0].check_mask.block[3].um_I.ena ,
    \top_I.branch[0].check_mask.block[2].um_I.ena ,
    \top_I.branch[0].check_mask.block[1].um_I.ena ,
    \top_I.branch[0].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[0].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[11].um_I.clk ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[10].um_I.clk ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[9].um_I.clk ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[8].um_I.clk ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[7].um_I.clk ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[6].um_I.clk ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[5].um_I.clk ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[4].um_I.clk ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[3].um_I.clk ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[2].um_I.clk ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[1].um_I.clk ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[0].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[0].um_I.pg_ena }));
 tt_pg_1v5_ll_2 \top_I.branch[10].check_mask.block[0].um_I.block_10_0.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[10].check_mask.block[0].um_I.block_10_0.vdpwr ),
    .ctrl(\top_I.branch[10].check_mask.block[0].um_I.pg_ena ));
 tt_um_rejunity_vga_logo \top_I.branch[10].check_mask.block[0].um_I.block_10_0.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[10].check_mask.block[0].um_I.block_10_0.vdpwr ),
    .clk(\top_I.branch[10].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[10].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[10].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[10].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[10].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[10].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[10].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[10].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[0] }));
 tt_pg_1v5_ll_2 \top_I.branch[10].check_mask.block[2].um_I.block_10_2.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[10].check_mask.block[2].um_I.block_10_2.vdpwr ),
    .ctrl(\top_I.branch[10].check_mask.block[2].um_I.pg_ena ));
 tt_um_rebeccargb_vga_pride \top_I.branch[10].check_mask.block[2].um_I.block_10_2.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[10].check_mask.block[2].um_I.block_10_2.vdpwr ),
    .clk(\top_I.branch[10].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[10].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[10].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[10].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[10].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[10].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[10].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[10].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[0] }));
 tt_mux \top_I.branch[10].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[10].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[10].check_mask.l_addr[1] ),
    .addr({\top_I.branch[10].check_mask.l_addr[1] ,
    \top_I.branch[10].check_mask.l_addr[0] ,
    \top_I.branch[10].check_mask.l_addr[1] ,
    \top_I.branch[10].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[10].check_mask.block[11].um_I.ena ,
    \top_I.branch[10].check_mask.block[10].um_I.ena ,
    \top_I.branch[10].check_mask.block[9].um_I.ena ,
    \top_I.branch[10].check_mask.block[8].um_I.ena ,
    \top_I.branch[10].check_mask.block[7].um_I.ena ,
    \top_I.branch[10].check_mask.block[6].um_I.ena ,
    \top_I.branch[10].check_mask.block[5].um_I.ena ,
    \top_I.branch[10].check_mask.block[4].um_I.ena ,
    \top_I.branch[10].check_mask.block[3].um_I.ena ,
    \top_I.branch[10].check_mask.block[2].um_I.ena ,
    \top_I.branch[10].check_mask.block[1].um_I.ena ,
    \top_I.branch[10].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[10].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[11].um_I.clk ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[10].um_I.clk ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[9].um_I.clk ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[8].um_I.clk ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[7].um_I.clk ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[6].um_I.clk ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[5].um_I.clk ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[4].um_I.clk ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[3].um_I.clk ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[2].um_I.clk ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[1].um_I.clk ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[10].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[13].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[13].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[13].check_mask.l_addr[0] ),
    .addr({\top_I.branch[13].check_mask.l_addr[0] ,
    \top_I.branch[13].check_mask.l_addr[1] ,
    \top_I.branch[13].check_mask.l_addr[1] ,
    \top_I.branch[13].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[13].check_mask.block[11].um_I.ena ,
    \top_I.branch[13].check_mask.block[10].um_I.ena ,
    \top_I.branch[13].check_mask.block[9].um_I.ena ,
    \top_I.branch[13].check_mask.block[8].um_I.ena ,
    \top_I.branch[13].check_mask.block[7].um_I.ena ,
    \top_I.branch[13].check_mask.block[6].um_I.ena ,
    \top_I.branch[13].check_mask.block[5].um_I.ena ,
    \top_I.branch[13].check_mask.block[4].um_I.ena ,
    \top_I.branch[13].check_mask.block[3].um_I.ena ,
    \top_I.branch[13].check_mask.block[2].um_I.ena ,
    \top_I.branch[13].check_mask.block[1].um_I.ena ,
    \top_I.branch[13].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[13].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[11].um_I.clk ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[10].um_I.clk ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[9].um_I.clk ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[8].um_I.clk ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[7].um_I.clk ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[6].um_I.clk ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[5].um_I.clk ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[4].um_I.clk ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[3].um_I.clk ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[2].um_I.clk ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[1].um_I.clk ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[13].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[14].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[14].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[14].check_mask.l_addr[3] ),
    .addr({\top_I.branch[14].check_mask.l_addr[3] ,
    \top_I.branch[14].check_mask.l_addr[0] ,
    \top_I.branch[14].check_mask.l_addr[0] ,
    \top_I.branch[14].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[14].check_mask.block[11].um_I.ena ,
    \top_I.branch[14].check_mask.block[10].um_I.ena ,
    \top_I.branch[14].check_mask.block[9].um_I.ena ,
    \top_I.branch[14].check_mask.block[8].um_I.ena ,
    \top_I.branch[14].check_mask.block[7].um_I.ena ,
    \top_I.branch[14].check_mask.block[6].um_I.ena ,
    \top_I.branch[14].check_mask.block[5].um_I.ena ,
    \top_I.branch[14].check_mask.block[4].um_I.ena ,
    \top_I.branch[14].check_mask.block[3].um_I.ena ,
    \top_I.branch[14].check_mask.block[2].um_I.ena ,
    \top_I.branch[14].check_mask.block[1].um_I.ena ,
    \top_I.branch[14].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[14].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[11].um_I.clk ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[10].um_I.clk ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[9].um_I.clk ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[8].um_I.clk ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[7].um_I.clk ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[6].um_I.clk ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[5].um_I.clk ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[4].um_I.clk ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[3].um_I.clk ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[2].um_I.clk ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[1].um_I.clk ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[14].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[15].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[15].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[15].check_mask.l_addr[3] ),
    .addr({\top_I.branch[15].check_mask.l_addr[3] ,
    \top_I.branch[15].check_mask.l_addr[0] ,
    \top_I.branch[15].check_mask.l_addr[0] ,
    \top_I.branch[15].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[15].check_mask.block[11].um_I.ena ,
    \top_I.branch[15].check_mask.block[10].um_I.ena ,
    \top_I.branch[15].check_mask.block[9].um_I.ena ,
    \top_I.branch[15].check_mask.block[8].um_I.ena ,
    \top_I.branch[15].check_mask.block[7].um_I.ena ,
    \top_I.branch[15].check_mask.block[6].um_I.ena ,
    \top_I.branch[15].check_mask.block[5].um_I.ena ,
    \top_I.branch[15].check_mask.block[4].um_I.ena ,
    \top_I.branch[15].check_mask.block[3].um_I.ena ,
    \top_I.branch[15].check_mask.block[2].um_I.ena ,
    \top_I.branch[15].check_mask.block[1].um_I.ena ,
    \top_I.branch[15].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[15].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[11].um_I.clk ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[10].um_I.clk ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[9].um_I.clk ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[8].um_I.clk ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[7].um_I.clk ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[6].um_I.clk ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[5].um_I.clk ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[4].um_I.clk ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[3].um_I.clk ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[2].um_I.clk ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[1].um_I.clk ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[15].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[0].um_I.pg_ena }));
 tt_pg_1v5_ll_1 \top_I.branch[16].check_mask.block[11].um_I.block_16_11.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[16].check_mask.block[11].um_I.block_16_11.vdpwr ),
    .ctrl(\top_I.branch[16].check_mask.block[11].um_I.pg_ena ));
 tt_um_rebeccargb_universal_decoder \top_I.branch[16].check_mask.block[11].um_I.block_16_11.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[16].check_mask.block[11].um_I.block_16_11.vdpwr ),
    .clk(\top_I.branch[16].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[0] }));
 tt_pg_1v5_ll_1 \top_I.branch[16].check_mask.block[1].um_I.block_16_1.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[16].check_mask.block[1].um_I.block_16_1.vdpwr ),
    .ctrl(\top_I.branch[16].check_mask.block[1].um_I.pg_ena ));
 tt_um_aksp_mbist_mbisr \top_I.branch[16].check_mask.block[1].um_I.block_16_1.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[16].check_mask.block[1].um_I.block_16_1.vdpwr ),
    .clk(\top_I.branch[16].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[0] }));
 tt_pg_1v5_ll_1 \top_I.branch[16].check_mask.block[3].um_I.block_16_3.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[16].check_mask.block[3].um_I.block_16_3.vdpwr ),
    .ctrl(\top_I.branch[16].check_mask.block[3].um_I.pg_ena ));
 tt_um_silicon_art \top_I.branch[16].check_mask.block[3].um_I.block_16_3.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[16].check_mask.block[3].um_I.block_16_3.vdpwr ),
    .clk(\top_I.branch[16].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[0] }));
 tt_pg_1v5_ll_1 \top_I.branch[16].check_mask.block[5].um_I.block_16_5.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[16].check_mask.block[5].um_I.block_16_5.vdpwr ),
    .ctrl(\top_I.branch[16].check_mask.block[5].um_I.pg_ena ));
 tt_um_urish_simon \top_I.branch[16].check_mask.block[5].um_I.block_16_5.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[16].check_mask.block[5].um_I.block_16_5.vdpwr ),
    .clk(\top_I.branch[16].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[0] }));
 tt_pg_1v5_ll_1 \top_I.branch[16].check_mask.block[7].um_I.block_16_7.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[16].check_mask.block[7].um_I.block_16_7.vdpwr ),
    .ctrl(\top_I.branch[16].check_mask.block[7].um_I.pg_ena ));
 tt_um_rebeccargb_intercal_alu \top_I.branch[16].check_mask.block[7].um_I.block_16_7.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[16].check_mask.block[7].um_I.block_16_7.vdpwr ),
    .clk(\top_I.branch[16].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[0] }));
 tt_pg_1v5_ll_1 \top_I.branch[16].check_mask.block[9].um_I.block_16_9.tt_pg_vdd_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .GPWR(\top_I.branch[16].check_mask.block[9].um_I.block_16_9.vdpwr ),
    .ctrl(\top_I.branch[16].check_mask.block[9].um_I.pg_ena ));
 tt_um_rebeccargb_hardware_utf8 \top_I.branch[16].check_mask.block[9].um_I.block_16_9.tt_um_I  (.VGND(vgnd),
    .VPWR(\top_I.branch[16].check_mask.block[9].um_I.block_16_9.vdpwr ),
    .clk(\top_I.branch[16].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[16].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[16].check_mask.l_addr[3] ),
    .k_zero(\top_I.branch[16].check_mask.l_addr[0] ),
    .addr({\top_I.branch[16].check_mask.l_addr[3] ,
    \top_I.branch[16].check_mask.l_addr[0] ,
    \top_I.branch[16].check_mask.l_addr[0] ,
    \top_I.branch[16].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[16].check_mask.block[11].um_I.ena ,
    \top_I.branch[16].check_mask.block[10].um_I.ena ,
    \top_I.branch[16].check_mask.block[9].um_I.ena ,
    \top_I.branch[16].check_mask.block[8].um_I.ena ,
    \top_I.branch[16].check_mask.block[7].um_I.ena ,
    \top_I.branch[16].check_mask.block[6].um_I.ena ,
    \top_I.branch[16].check_mask.block[5].um_I.ena ,
    \top_I.branch[16].check_mask.block[4].um_I.ena ,
    \top_I.branch[16].check_mask.block[3].um_I.ena ,
    \top_I.branch[16].check_mask.block[2].um_I.ena ,
    \top_I.branch[16].check_mask.block[1].um_I.ena ,
    \top_I.branch[16].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[16].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[11].um_I.clk ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[10].um_I.clk ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[9].um_I.clk ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[8].um_I.clk ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[7].um_I.clk ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[6].um_I.clk ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[5].um_I.clk ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[4].um_I.clk ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[3].um_I.clk ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[2].um_I.clk ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[1].um_I.clk ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[16].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[16].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[17].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[17].check_mask.l_addr[3] ),
    .k_zero(\top_I.branch[17].check_mask.l_addr[0] ),
    .addr({\top_I.branch[17].check_mask.l_addr[3] ,
    \top_I.branch[17].check_mask.l_addr[0] ,
    \top_I.branch[17].check_mask.l_addr[0] ,
    \top_I.branch[17].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[17].check_mask.block[11].um_I.ena ,
    \top_I.branch[17].check_mask.block[10].um_I.ena ,
    \top_I.branch[17].check_mask.block[9].um_I.ena ,
    \top_I.branch[17].check_mask.block[8].um_I.ena ,
    \top_I.branch[17].check_mask.block[7].um_I.ena ,
    \top_I.branch[17].check_mask.block[6].um_I.ena ,
    \top_I.branch[17].check_mask.block[5].um_I.ena ,
    \top_I.branch[17].check_mask.block[4].um_I.ena ,
    \top_I.branch[17].check_mask.block[3].um_I.ena ,
    \top_I.branch[17].check_mask.block[2].um_I.ena ,
    \top_I.branch[17].check_mask.block[1].um_I.ena ,
    \top_I.branch[17].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[17].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[11].um_I.clk ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[10].um_I.clk ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[9].um_I.clk ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[8].um_I.clk ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[7].um_I.clk ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[6].um_I.clk ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[5].um_I.clk ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[4].um_I.clk ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[3].um_I.clk ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[2].um_I.clk ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[1].um_I.clk ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[17].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[18].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[18].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[18].check_mask.l_addr[1] ),
    .addr({\top_I.branch[18].check_mask.l_addr[0] ,
    \top_I.branch[18].check_mask.l_addr[1] ,
    \top_I.branch[18].check_mask.l_addr[1] ,
    \top_I.branch[18].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[18].check_mask.block[11].um_I.ena ,
    \top_I.branch[18].check_mask.block[10].um_I.ena ,
    \top_I.branch[18].check_mask.block[9].um_I.ena ,
    \top_I.branch[18].check_mask.block[8].um_I.ena ,
    \top_I.branch[18].check_mask.block[7].um_I.ena ,
    \top_I.branch[18].check_mask.block[6].um_I.ena ,
    \top_I.branch[18].check_mask.block[5].um_I.ena ,
    \top_I.branch[18].check_mask.block[4].um_I.ena ,
    \top_I.branch[18].check_mask.block[3].um_I.ena ,
    \top_I.branch[18].check_mask.block[2].um_I.ena ,
    \top_I.branch[18].check_mask.block[1].um_I.ena ,
    \top_I.branch[18].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[18].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[11].um_I.clk ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[10].um_I.clk ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[9].um_I.clk ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[8].um_I.clk ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[7].um_I.clk ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[6].um_I.clk ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[5].um_I.clk ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[4].um_I.clk ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[3].um_I.clk ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[2].um_I.clk ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[1].um_I.clk ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[18].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[19].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[19].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[19].check_mask.l_addr[1] ),
    .addr({\top_I.branch[19].check_mask.l_addr[0] ,
    \top_I.branch[19].check_mask.l_addr[1] ,
    \top_I.branch[19].check_mask.l_addr[1] ,
    \top_I.branch[19].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[19].check_mask.block[11].um_I.ena ,
    \top_I.branch[19].check_mask.block[10].um_I.ena ,
    \top_I.branch[19].check_mask.block[9].um_I.ena ,
    \top_I.branch[19].check_mask.block[8].um_I.ena ,
    \top_I.branch[19].check_mask.block[7].um_I.ena ,
    \top_I.branch[19].check_mask.block[6].um_I.ena ,
    \top_I.branch[19].check_mask.block[5].um_I.ena ,
    \top_I.branch[19].check_mask.block[4].um_I.ena ,
    \top_I.branch[19].check_mask.block[3].um_I.ena ,
    \top_I.branch[19].check_mask.block[2].um_I.ena ,
    \top_I.branch[19].check_mask.block[1].um_I.ena ,
    \top_I.branch[19].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[19].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[11].um_I.clk ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[10].um_I.clk ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[9].um_I.clk ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[8].um_I.clk ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[7].um_I.clk ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[6].um_I.clk ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[5].um_I.clk ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[4].um_I.clk ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[3].um_I.clk ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[2].um_I.clk ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[1].um_I.clk ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[19].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[1].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[1].check_mask.l_k_one ),
    .k_zero(\top_I.branch[1].check_mask.l_addr[0] ),
    .addr({\top_I.branch[1].check_mask.l_addr[0] ,
    \top_I.branch[1].check_mask.l_addr[0] ,
    \top_I.branch[1].check_mask.l_addr[0] ,
    \top_I.branch[1].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[1].check_mask.block[11].um_I.ena ,
    \top_I.branch[1].check_mask.block[10].um_I.ena ,
    \top_I.branch[1].check_mask.block[9].um_I.ena ,
    \top_I.branch[1].check_mask.block[8].um_I.ena ,
    \top_I.branch[1].check_mask.block[7].um_I.ena ,
    \top_I.branch[1].check_mask.block[6].um_I.ena ,
    \top_I.branch[1].check_mask.block[5].um_I.ena ,
    \top_I.branch[1].check_mask.block[4].um_I.ena ,
    \top_I.branch[1].check_mask.block[3].um_I.ena ,
    \top_I.branch[1].check_mask.block[2].um_I.ena ,
    \top_I.branch[1].check_mask.block[1].um_I.ena ,
    \top_I.branch[1].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[1].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[11].um_I.clk ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[10].um_I.clk ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[9].um_I.clk ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[8].um_I.clk ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[7].um_I.clk ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[6].um_I.clk ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[5].um_I.clk ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[4].um_I.clk ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[3].um_I.clk ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[2].um_I.clk ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[1].um_I.clk ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[1].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[2].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[2].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[2].check_mask.l_addr[1] ),
    .addr({\top_I.branch[2].check_mask.l_addr[1] ,
    \top_I.branch[2].check_mask.l_addr[1] ,
    \top_I.branch[2].check_mask.l_addr[1] ,
    \top_I.branch[2].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[2].check_mask.block[11].um_I.ena ,
    \top_I.branch[2].check_mask.block[10].um_I.ena ,
    \top_I.branch[2].check_mask.block[9].um_I.ena ,
    \top_I.branch[2].check_mask.block[8].um_I.ena ,
    \top_I.branch[2].check_mask.block[7].um_I.ena ,
    \top_I.branch[2].check_mask.block[6].um_I.ena ,
    \top_I.branch[2].check_mask.block[5].um_I.ena ,
    \top_I.branch[2].check_mask.block[4].um_I.ena ,
    \top_I.branch[2].check_mask.block[3].um_I.ena ,
    \top_I.branch[2].check_mask.block[2].um_I.ena ,
    \top_I.branch[2].check_mask.block[1].um_I.ena ,
    \top_I.branch[2].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[2].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[11].um_I.clk ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[10].um_I.clk ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[9].um_I.clk ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[8].um_I.clk ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[7].um_I.clk ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[6].um_I.clk ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[5].um_I.clk ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[4].um_I.clk ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[3].um_I.clk ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[2].um_I.clk ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[1].um_I.clk ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[2].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[3].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[3].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[3].check_mask.l_addr[1] ),
    .addr({\top_I.branch[3].check_mask.l_addr[1] ,
    \top_I.branch[3].check_mask.l_addr[1] ,
    \top_I.branch[3].check_mask.l_addr[1] ,
    \top_I.branch[3].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[3].check_mask.block[11].um_I.ena ,
    \top_I.branch[3].check_mask.block[10].um_I.ena ,
    \top_I.branch[3].check_mask.block[9].um_I.ena ,
    \top_I.branch[3].check_mask.block[8].um_I.ena ,
    \top_I.branch[3].check_mask.block[7].um_I.ena ,
    \top_I.branch[3].check_mask.block[6].um_I.ena ,
    \top_I.branch[3].check_mask.block[5].um_I.ena ,
    \top_I.branch[3].check_mask.block[4].um_I.ena ,
    \top_I.branch[3].check_mask.block[3].um_I.ena ,
    \top_I.branch[3].check_mask.block[2].um_I.ena ,
    \top_I.branch[3].check_mask.block[1].um_I.ena ,
    \top_I.branch[3].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[3].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[11].um_I.clk ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[10].um_I.clk ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[9].um_I.clk ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[8].um_I.clk ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[7].um_I.clk ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[6].um_I.clk ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[5].um_I.clk ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[4].um_I.clk ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[3].um_I.clk ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[2].um_I.clk ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[1].um_I.clk ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[3].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[4].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[4].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[4].check_mask.l_addr[0] ),
    .addr({\top_I.branch[4].check_mask.l_addr[0] ,
    \top_I.branch[4].check_mask.l_addr[0] ,
    \top_I.branch[4].check_mask.l_addr[1] ,
    \top_I.branch[4].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[4].check_mask.block[11].um_I.ena ,
    \top_I.branch[4].check_mask.block[10].um_I.ena ,
    \top_I.branch[4].check_mask.block[9].um_I.ena ,
    \top_I.branch[4].check_mask.block[8].um_I.ena ,
    \top_I.branch[4].check_mask.block[7].um_I.ena ,
    \top_I.branch[4].check_mask.block[6].um_I.ena ,
    \top_I.branch[4].check_mask.block[5].um_I.ena ,
    \top_I.branch[4].check_mask.block[4].um_I.ena ,
    \top_I.branch[4].check_mask.block[3].um_I.ena ,
    \top_I.branch[4].check_mask.block[2].um_I.ena ,
    \top_I.branch[4].check_mask.block[1].um_I.ena ,
    \top_I.branch[4].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[4].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[11].um_I.clk ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[10].um_I.clk ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[9].um_I.clk ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[8].um_I.clk ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[7].um_I.clk ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[6].um_I.clk ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[5].um_I.clk ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[4].um_I.clk ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[3].um_I.clk ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[2].um_I.clk ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[1].um_I.clk ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[4].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[5].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[5].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[5].check_mask.l_addr[0] ),
    .addr({\top_I.branch[5].check_mask.l_addr[0] ,
    \top_I.branch[5].check_mask.l_addr[0] ,
    \top_I.branch[5].check_mask.l_addr[1] ,
    \top_I.branch[5].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[5].check_mask.block[11].um_I.ena ,
    \top_I.branch[5].check_mask.block[10].um_I.ena ,
    \top_I.branch[5].check_mask.block[9].um_I.ena ,
    \top_I.branch[5].check_mask.block[8].um_I.ena ,
    \top_I.branch[5].check_mask.block[7].um_I.ena ,
    \top_I.branch[5].check_mask.block[6].um_I.ena ,
    \top_I.branch[5].check_mask.block[5].um_I.ena ,
    \top_I.branch[5].check_mask.block[4].um_I.ena ,
    \top_I.branch[5].check_mask.block[3].um_I.ena ,
    \top_I.branch[5].check_mask.block[2].um_I.ena ,
    \top_I.branch[5].check_mask.block[1].um_I.ena ,
    \top_I.branch[5].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[5].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[11].um_I.clk ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[10].um_I.clk ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[9].um_I.clk ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[8].um_I.clk ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[7].um_I.clk ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[6].um_I.clk ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[5].um_I.clk ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[4].um_I.clk ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[3].um_I.clk ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[2].um_I.clk ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[1].um_I.clk ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[5].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[7].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[7].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[7].check_mask.l_addr[2] ),
    .addr({\top_I.branch[7].check_mask.l_addr[2] ,
    \top_I.branch[7].check_mask.l_addr[2] ,
    \top_I.branch[7].check_mask.l_addr[0] ,
    \top_I.branch[7].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[7].check_mask.block[11].um_I.ena ,
    \top_I.branch[7].check_mask.block[10].um_I.ena ,
    \top_I.branch[7].check_mask.block[9].um_I.ena ,
    \top_I.branch[7].check_mask.block[8].um_I.ena ,
    \top_I.branch[7].check_mask.block[7].um_I.ena ,
    \top_I.branch[7].check_mask.block[6].um_I.ena ,
    \top_I.branch[7].check_mask.block[5].um_I.ena ,
    \top_I.branch[7].check_mask.block[4].um_I.ena ,
    \top_I.branch[7].check_mask.block[3].um_I.ena ,
    \top_I.branch[7].check_mask.block[2].um_I.ena ,
    \top_I.branch[7].check_mask.block[1].um_I.ena ,
    \top_I.branch[7].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[7].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[11].um_I.clk ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[10].um_I.clk ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[9].um_I.clk ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[8].um_I.clk ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[7].um_I.clk ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[6].um_I.clk ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[5].um_I.clk ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[4].um_I.clk ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[3].um_I.clk ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[2].um_I.clk ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[1].um_I.clk ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[7].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[8].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[8].check_mask.l_addr[2] ),
    .k_zero(\top_I.branch[8].check_mask.l_addr[0] ),
    .addr({\top_I.branch[8].check_mask.l_addr[0] ,
    \top_I.branch[8].check_mask.l_addr[2] ,
    \top_I.branch[8].check_mask.l_addr[0] ,
    \top_I.branch[8].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[8].check_mask.block[11].um_I.ena ,
    \top_I.branch[8].check_mask.block[10].um_I.ena ,
    \top_I.branch[8].check_mask.block[9].um_I.ena ,
    \top_I.branch[8].check_mask.block[8].um_I.ena ,
    \top_I.branch[8].check_mask.block[7].um_I.ena ,
    \top_I.branch[8].check_mask.block[6].um_I.ena ,
    \top_I.branch[8].check_mask.block[5].um_I.ena ,
    \top_I.branch[8].check_mask.block[4].um_I.ena ,
    \top_I.branch[8].check_mask.block[3].um_I.ena ,
    \top_I.branch[8].check_mask.block[2].um_I.ena ,
    \top_I.branch[8].check_mask.block[1].um_I.ena ,
    \top_I.branch[8].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[8].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[11].um_I.clk ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[10].um_I.clk ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[9].um_I.clk ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[8].um_I.clk ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[7].um_I.clk ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[6].um_I.clk ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[5].um_I.clk ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[4].um_I.clk ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[3].um_I.clk ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[2].um_I.clk ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[1].um_I.clk ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[8].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[0].um_I.pg_ena }));
 tt_mux \top_I.branch[9].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[9].check_mask.l_addr[2] ),
    .k_zero(\top_I.branch[9].check_mask.l_addr[0] ),
    .addr({\top_I.branch[9].check_mask.l_addr[0] ,
    \top_I.branch[9].check_mask.l_addr[2] ,
    \top_I.branch[9].check_mask.l_addr[0] ,
    \top_I.branch[9].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[9].check_mask.block[11].um_I.ena ,
    \top_I.branch[9].check_mask.block[10].um_I.ena ,
    \top_I.branch[9].check_mask.block[9].um_I.ena ,
    \top_I.branch[9].check_mask.block[8].um_I.ena ,
    \top_I.branch[9].check_mask.block[7].um_I.ena ,
    \top_I.branch[9].check_mask.block[6].um_I.ena ,
    \top_I.branch[9].check_mask.block[5].um_I.ena ,
    \top_I.branch[9].check_mask.block[4].um_I.ena ,
    \top_I.branch[9].check_mask.block[3].um_I.ena ,
    \top_I.branch[9].check_mask.block[2].um_I.ena ,
    \top_I.branch[9].check_mask.block[1].um_I.ena ,
    \top_I.branch[9].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[9].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[11].um_I.clk ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[10].um_I.clk ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[9].um_I.clk ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[8].um_I.clk ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[7].um_I.clk ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[6].um_I.clk ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[5].um_I.clk ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[4].um_I.clk ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[3].um_I.clk ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[2].um_I.clk ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[1].um_I.clk ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[9].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[0].um_I.pg_ena }));
 tt_ctrl \top_I.ctrl_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .ctrl_ena(\gpio[0].gpio_I.pad_in ),
    .ctrl_sel_inc(\gpio[1].gpio_I.pad_in ),
    .ctrl_sel_rst_n(\gpio[2].gpio_I.pad_in ),
    .k_one(\gpio[0].gpio_I.pad_oe ),
    .k_zero(\gpio[18].gpio_I.pad_oe ),
    .pad_ui_in({\gpio[47].gpio_I.pad_in ,
    \gpio[46].gpio_I.pad_in ,
    \gpio[45].gpio_I.pad_in ,
    \gpio[44].gpio_I.pad_in ,
    \gpio[43].gpio_I.pad_in ,
    \gpio[42].gpio_I.pad_in ,
    \gpio[41].gpio_I.pad_in ,
    \gpio[40].gpio_I.pad_in ,
    \gpio[48].gpio_I.pad_in ,
    \gpio[49].gpio_I.pad_in }),
    .pad_uio_in({\gpio[39].gpio_I.pad_in ,
    \gpio[38].gpio_I.pad_in ,
    \gpio[37].gpio_I.pad_in ,
    \gpio[36].gpio_I.pad_in ,
    \gpio[35].gpio_I.pad_in ,
    \gpio[34].gpio_I.pad_in ,
    \gpio[33].gpio_I.pad_in ,
    \gpio[32].gpio_I.pad_in }),
    .pad_uio_oex({\gpio[39].gpio_I.pad_oe ,
    \gpio[38].gpio_I.pad_oe ,
    \gpio[37].gpio_I.pad_oe ,
    \gpio[36].gpio_I.pad_oe ,
    \gpio[35].gpio_I.pad_oe ,
    \gpio[34].gpio_I.pad_oe ,
    \gpio[33].gpio_I.pad_oe ,
    \gpio[32].gpio_I.pad_oe }),
    .pad_uio_out({\gpio[39].gpio_I.pad_out ,
    \gpio[38].gpio_I.pad_out ,
    \gpio[37].gpio_I.pad_out ,
    \gpio[36].gpio_I.pad_out ,
    \gpio[35].gpio_I.pad_out ,
    \gpio[34].gpio_I.pad_out ,
    \gpio[33].gpio_I.pad_out ,
    \gpio[32].gpio_I.pad_out }),
    .pad_uo_out({\gpio[15].gpio_I.pad_out ,
    \gpio[14].gpio_I.pad_out ,
    \gpio[13].gpio_I.pad_out ,
    \gpio[12].gpio_I.pad_out ,
    \gpio[11].gpio_I.pad_out ,
    \gpio[10].gpio_I.pad_out ,
    \gpio[9].gpio_I.pad_out ,
    \gpio[8].gpio_I.pad_out }),
    .spine_bot_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_bot_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .spine_top_iw({\top_I.branch[13].check_mask.l_spine_iw[29] ,
    \top_I.branch[13].check_mask.l_spine_iw[28] ,
    \top_I.branch[13].check_mask.l_spine_iw[27] ,
    \top_I.branch[13].check_mask.l_spine_iw[26] ,
    \top_I.branch[13].check_mask.l_spine_iw[25] ,
    \top_I.branch[13].check_mask.l_spine_iw[24] ,
    \top_I.branch[13].check_mask.l_spine_iw[23] ,
    \top_I.branch[13].check_mask.l_spine_iw[22] ,
    \top_I.branch[13].check_mask.l_spine_iw[21] ,
    \top_I.branch[13].check_mask.l_spine_iw[20] ,
    \top_I.branch[13].check_mask.l_spine_iw[19] ,
    \top_I.branch[13].check_mask.l_spine_iw[18] ,
    \top_I.branch[13].check_mask.l_spine_iw[17] ,
    \top_I.branch[13].check_mask.l_spine_iw[16] ,
    \top_I.branch[13].check_mask.l_spine_iw[15] ,
    \top_I.branch[13].check_mask.l_spine_iw[14] ,
    \top_I.branch[13].check_mask.l_spine_iw[13] ,
    \top_I.branch[13].check_mask.l_spine_iw[12] ,
    \top_I.branch[13].check_mask.l_spine_iw[11] ,
    \top_I.branch[13].check_mask.l_spine_iw[10] ,
    \top_I.branch[13].check_mask.l_spine_iw[9] ,
    \top_I.branch[13].check_mask.l_spine_iw[8] ,
    \top_I.branch[13].check_mask.l_spine_iw[7] ,
    \top_I.branch[13].check_mask.l_spine_iw[6] ,
    \top_I.branch[13].check_mask.l_spine_iw[5] ,
    \top_I.branch[13].check_mask.l_spine_iw[4] ,
    \top_I.branch[13].check_mask.l_spine_iw[3] ,
    \top_I.branch[13].check_mask.l_spine_iw[2] ,
    \top_I.branch[13].check_mask.l_spine_iw[1] ,
    \top_I.branch[13].check_mask.l_spine_iw[0] }),
    .spine_top_ow({\top_I.branch[13].check_mask.l_spine_ow[25] ,
    \top_I.branch[13].check_mask.l_spine_ow[24] ,
    \top_I.branch[13].check_mask.l_spine_ow[23] ,
    \top_I.branch[13].check_mask.l_spine_ow[22] ,
    \top_I.branch[13].check_mask.l_spine_ow[21] ,
    \top_I.branch[13].check_mask.l_spine_ow[20] ,
    \top_I.branch[13].check_mask.l_spine_ow[19] ,
    \top_I.branch[13].check_mask.l_spine_ow[18] ,
    \top_I.branch[13].check_mask.l_spine_ow[17] ,
    \top_I.branch[13].check_mask.l_spine_ow[16] ,
    \top_I.branch[13].check_mask.l_spine_ow[15] ,
    \top_I.branch[13].check_mask.l_spine_ow[14] ,
    \top_I.branch[13].check_mask.l_spine_ow[13] ,
    \top_I.branch[13].check_mask.l_spine_ow[12] ,
    \top_I.branch[13].check_mask.l_spine_ow[11] ,
    \top_I.branch[13].check_mask.l_spine_ow[10] ,
    \top_I.branch[13].check_mask.l_spine_ow[9] ,
    \top_I.branch[13].check_mask.l_spine_ow[8] ,
    \top_I.branch[13].check_mask.l_spine_ow[7] ,
    \top_I.branch[13].check_mask.l_spine_ow[6] ,
    \top_I.branch[13].check_mask.l_spine_ow[5] ,
    \top_I.branch[13].check_mask.l_spine_ow[4] ,
    \top_I.branch[13].check_mask.l_spine_ow[3] ,
    \top_I.branch[13].check_mask.l_spine_ow[2] ,
    \top_I.branch[13].check_mask.l_spine_ow[1] ,
    \top_I.branch[13].check_mask.l_spine_ow[0] }));
 tt_logo_bottom \top_I.logo_bottom_I  ();
 tt_logo_corner \top_I.logo_corner_I  ();
 tt_logo_top \top_I.logo_top_I  ();
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_0_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_0_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_1_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_1_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_1_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_1_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_2_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_2_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_2_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_2_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_3_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_3_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_3_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_3_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_4_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_4_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_4_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_4_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_5_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_5_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_5_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_5_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_6_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_6_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_6_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_6_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_7_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_7_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_7_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_7_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_8_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_8_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_8_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_8_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_9_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_9_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_9_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_9_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_10_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_10_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_10_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_10_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_11_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_11_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_11_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_11_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_12_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_12_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_12_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_12_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_13_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_13_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_13_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_13_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_14_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_14_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_14_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_14_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_15_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_15_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_15_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_NORTH_15_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_16_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_16_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_0_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_0_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_1_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_1_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_1_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_1_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_2_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_2_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_2_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_2_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_3_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_3_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_3_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_3_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_4_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_4_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_4_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_4_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_5_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_5_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_5_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_5_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_6_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_6_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_6_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_6_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_7_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_7_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_7_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_7_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_8_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_8_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_8_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_8_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_9_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_9_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_9_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_9_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_10_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_10_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_10_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_10_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_11_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_11_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_11_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_11_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_12_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_12_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_12_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_12_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_13_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_13_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_13_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_13_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_14_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_14_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_14_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_14_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_15_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_15_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_15_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_SOUTH_15_102 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_16_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_16_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_0_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_0_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_1_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_1_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_1_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_1_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_1_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_1_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_2_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_2_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_2_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_2_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_2_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_2_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_3_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_3_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_3_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_3_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_3_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_3_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_4_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_4_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_4_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_4_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_4_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_4_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_5_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_5_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_5_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_5_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_5_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_5_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_6_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_6_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_6_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_6_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_6_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_6_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_7_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_7_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_7_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_7_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_7_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_7_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_8_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_8_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_8_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_8_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_8_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_8_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_9_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_9_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_9_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_9_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_9_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_9_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_10_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_10_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_10_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_10_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_10_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_10_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_11_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_11_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_11_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_11_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_11_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_11_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_12_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_12_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_12_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_12_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_12_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_12_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_13_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_13_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_13_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_13_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_13_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_13_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_14_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_14_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_14_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_14_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_14_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_14_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_15_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_15_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_15_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_15_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_15_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_15_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_16_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_16_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_0_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_0_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_1_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_1_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_1_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_1_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_1_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_1_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_2_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_2_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_2_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_2_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_2_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_2_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_3_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_3_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_3_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_3_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_3_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_3_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_4_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_4_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_4_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_4_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_4_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_4_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_5_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_5_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_5_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_5_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_5_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_5_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_6_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_6_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_6_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_6_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_6_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_6_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_7_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_7_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_7_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_7_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_7_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_7_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_8_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_8_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_8_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_8_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_8_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_8_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_9_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_9_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_9_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_9_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_9_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_9_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_10_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_10_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_10_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_10_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_10_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_10_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_11_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_11_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_11_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_11_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_11_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_11_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_12_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_12_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_12_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_12_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_12_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_12_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_13_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_13_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_13_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_13_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_13_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_13_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_14_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_14_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_14_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_14_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_14_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_14_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_15_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_15_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_15_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_15_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_15_170 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_15_190 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_16_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_16_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 bondpad_70x70 \IO_BOND_gpio[0].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[0]));
 bondpad_70x70 \IO_BOND_gpio[10].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[10]));
 bondpad_70x70 \IO_BOND_gpio[11].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[11]));
 bondpad_70x70 \IO_BOND_gpio[12].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[12]));
 bondpad_70x70 \IO_BOND_gpio[13].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[13]));
 bondpad_70x70 \IO_BOND_gpio[14].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[14]));
 bondpad_70x70 \IO_BOND_gpio[15].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[15]));
 bondpad_70x70 \IO_BOND_gpio[16].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[17].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[18].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[19].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[1].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[1]));
 bondpad_70x70 \IO_BOND_gpio[20].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[21].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[22].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[23].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[24].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[25].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[26].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[27].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[28].gpio_I.genblk1.pad_I  (.pad(vgnd));
 bondpad_70x70 \IO_BOND_gpio[29].gpio_I.genblk1.genblk1.pad_I  (.pad(vdpwr));
 bondpad_70x70 \IO_BOND_gpio[2].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[2]));
 bondpad_70x70 \IO_BOND_gpio[30].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[31].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[32].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[32]));
 bondpad_70x70 \IO_BOND_gpio[33].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[33]));
 bondpad_70x70 \IO_BOND_gpio[34].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[34]));
 bondpad_70x70 \IO_BOND_gpio[35].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[35]));
 bondpad_70x70 \IO_BOND_gpio[36].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[36]));
 bondpad_70x70 \IO_BOND_gpio[37].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[37]));
 bondpad_70x70 \IO_BOND_gpio[38].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[38]));
 bondpad_70x70 \IO_BOND_gpio[39].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[39]));
 bondpad_70x70 \IO_BOND_gpio[3].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[3]));
 bondpad_70x70 \IO_BOND_gpio[40].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[40]));
 bondpad_70x70 \IO_BOND_gpio[41].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[41]));
 bondpad_70x70 \IO_BOND_gpio[42].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[42]));
 bondpad_70x70 \IO_BOND_gpio[43].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[43]));
 bondpad_70x70 \IO_BOND_gpio[44].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[44]));
 bondpad_70x70 \IO_BOND_gpio[45].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[45]));
 bondpad_70x70 \IO_BOND_gpio[46].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[46]));
 bondpad_70x70 \IO_BOND_gpio[47].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[47]));
 bondpad_70x70 \IO_BOND_gpio[48].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[48]));
 bondpad_70x70 \IO_BOND_gpio[49].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[49]));
 bondpad_70x70 \IO_BOND_gpio[4].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[4]));
 bondpad_70x70 \IO_BOND_gpio[50].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[51].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[52].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[53].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[54].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[55].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[56].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[57].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[58].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[59].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[5].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[5]));
 bondpad_70x70 \IO_BOND_gpio[60].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[61].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[62].gpio_I.genblk1.pad_I  (.pad(vgnd));
 bondpad_70x70 \IO_BOND_gpio[63].gpio_I.genblk1.genblk1.pad_I  (.pad(vdpwr));
 bondpad_70x70 \IO_BOND_gpio[6].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[7].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[8].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[8]));
 bondpad_70x70 \IO_BOND_gpio[9].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk3.pad_I  (.pad(pad_raw[9]));
endmodule
